module GraphReader(
  input        clock,
  input        reset,
  input        io_valid_in,
  output       io_valid_out,
  input        io_flag_job,
  input  [2:0] io_job_big_bank_id,
  input  [9:0] io_job_big_cnt_x_end,
  input  [9:0] io_job_big_cnt_y_end,
  input  [9:0] io_job_big_cnt_ic_end,
  input  [9:0] io_job_big_cnt_loop_end,
  input  [9:0] io_job_big_begin_loop,
  input  [9:0] io_job_small_0_max_addr,
  input  [9:0] io_job_small_0_cnt_y_end,
  input  [9:0] io_job_small_0_cnt_ic_end,
  input  [9:0] io_job_small_0_cnt_loop_end,
  input  [9:0] io_job_small_0_begin_loop,
  input  [9:0] io_job_small_0_cnt_invalid_end,
  output [2:0] io_to_banks_addrs_0_bank_id,
  output [9:0] io_to_banks_addrs_1_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] gen_big_cnt_ic_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_big_cnt_ic_cend; // @[read.scala 26:22]
  reg [9:0] gen_big_cnt_x_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_big_cnt_x_cend; // @[read.scala 26:22]
  reg [9:0] gen_big_cnt_y_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_big_cnt_y_cend; // @[read.scala 26:22]
  reg [2:0] gen_big_bank_id; // @[read.scala 26:22]
  reg [9:0] gen_big_cnt_loop_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_big_cnt_loop_cend; // @[read.scala 26:22]
  reg  gen_big_cnt_ups_ccnt; // @[read.scala 26:22]
  reg  gen_big_flag_end; // @[read.scala 26:22]
  reg [9:0] gen_small_0_max_addr; // @[read.scala 26:22]
  reg [9:0] gen_small_0_now_addr; // @[read.scala 26:22]
  reg [9:0] gen_small_0_cnt_ic_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_small_0_cnt_ic_cend; // @[read.scala 26:22]
  reg [9:0] gen_small_0_cnt_y_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_small_0_cnt_y_cend; // @[read.scala 26:22]
  reg [9:0] gen_small_0_cnt_invalid_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_small_0_cnt_invalid_cend; // @[read.scala 26:22]
  reg  gen_small_0_cnt_ups_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_small_0_cnt_loop_ccnt; // @[read.scala 26:22]
  reg [9:0] gen_small_0_cnt_loop_cend; // @[read.scala 26:22]
  reg  gen_small_0_cnt_swap_ccnt; // @[read.scala 26:22]
  reg  gen_small_0_cnt_swap_cend; // @[read.scala 26:22]
  reg [9:0] gen_small_0_y_begin_addr; // @[read.scala 26:22]
  reg [9:0] gen_small_0_ic_begin_addr; // @[read.scala 26:22]
  reg  gen_small_0_start; // @[read.scala 26:22]
  wire  nxt = gen_big_cnt_ic_ccnt == gen_big_cnt_ic_cend; // @[utils.scala 17:20]
  wire [9:0] _gen_big_cnt_ic_ccnt_T_1 = gen_big_cnt_ic_ccnt + 10'h1; // @[utils.scala 18:35]
  wire  nxt_1 = gen_big_cnt_loop_ccnt == gen_big_cnt_loop_cend; // @[utils.scala 17:20]
  wire [9:0] _gen_big_cnt_loop_ccnt_T_1 = gen_big_cnt_loop_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_big_cnt_loop_ccnt_T_2 = nxt_1 ? 10'h0 : _gen_big_cnt_loop_ccnt_T_1; // @[utils.scala 18:20]
  wire  nxt_2 = gen_big_cnt_y_ccnt == gen_big_cnt_y_cend; // @[utils.scala 17:20]
  wire [9:0] _gen_big_cnt_y_ccnt_T_1 = gen_big_cnt_y_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_big_cnt_y_ccnt_T_2 = nxt_2 ? 10'h0 : _gen_big_cnt_y_ccnt_T_1; // @[utils.scala 18:20]
  wire  nxt_3 = ~gen_big_cnt_ups_ccnt; // @[utils.scala 17:20]
  wire  _gen_big_cnt_ups_ccnt_T_2 = nxt_3 ? 1'h0 : gen_big_cnt_ups_ccnt + 1'h1; // @[utils.scala 18:20]
  wire  nxt_4 = gen_big_cnt_x_ccnt == gen_big_cnt_x_cend; // @[utils.scala 17:20]
  wire [9:0] _gen_big_cnt_x_ccnt_T_1 = gen_big_cnt_x_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_big_cnt_x_ccnt_T_2 = nxt_4 ? 10'h0 : _gen_big_cnt_x_ccnt_T_1; // @[utils.scala 18:20]
  wire  _GEN_0 = nxt_4 | gen_big_flag_end; // @[gen_addr.scala 85:42 gen_addr.scala 86:38 read.scala 26:22]
  wire [9:0] _GEN_3 = nxt_3 ? _gen_big_cnt_x_ccnt_T_2 : gen_big_cnt_x_ccnt; // @[gen_addr.scala 84:40 utils.scala 18:14 read.scala 26:22]
  wire  _GEN_4 = nxt_3 ? _GEN_0 : gen_big_flag_end; // @[gen_addr.scala 84:40 read.scala 26:22]
  wire  _GEN_7 = nxt_2 ? _gen_big_cnt_ups_ccnt_T_2 : gen_big_cnt_ups_ccnt; // @[gen_addr.scala 83:34 utils.scala 18:14 read.scala 26:22]
  wire [9:0] _GEN_8 = nxt_2 ? _GEN_3 : gen_big_cnt_x_ccnt; // @[gen_addr.scala 83:34 read.scala 26:22]
  wire  _GEN_9 = nxt_2 ? _GEN_4 : gen_big_flag_end; // @[gen_addr.scala 83:34 read.scala 26:22]
  wire [9:0] _GEN_13 = nxt_1 ? _gen_big_cnt_y_ccnt_T_2 : gen_big_cnt_y_ccnt; // @[gen_addr.scala 82:33 utils.scala 18:14 read.scala 26:22]
  wire  _GEN_14 = nxt_1 ? _GEN_7 : gen_big_cnt_ups_ccnt; // @[gen_addr.scala 82:33 read.scala 26:22]
  wire [9:0] _GEN_15 = nxt_1 ? _GEN_8 : gen_big_cnt_x_ccnt; // @[gen_addr.scala 82:33 read.scala 26:22]
  wire  _GEN_16 = nxt_1 ? _GEN_9 : gen_big_flag_end; // @[gen_addr.scala 82:33 read.scala 26:22]
  wire  nxt_5 = gen_small_0_cnt_invalid_ccnt == gen_small_0_cnt_invalid_cend; // @[utils.scala 17:20]
  wire [9:0] _gen_small_0_cnt_invalid_ccnt_T_1 = gen_small_0_cnt_invalid_ccnt + 10'h1; // @[utils.scala 18:35]
  wire  nxt_6 = gen_small_0_cnt_ic_ccnt == gen_small_0_cnt_ic_cend; // @[utils.scala 17:20]
  wire [9:0] _gen_small_0_cnt_ic_ccnt_T_1 = gen_small_0_cnt_ic_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_small_0_cnt_ic_ccnt_T_2 = nxt_6 ? 10'h0 : _gen_small_0_cnt_ic_ccnt_T_1; // @[utils.scala 18:20]
  wire  nxt_7 = gen_small_0_cnt_loop_ccnt == gen_small_0_cnt_loop_cend; // @[utils.scala 17:20]
  wire [9:0] _gen_small_0_cnt_loop_ccnt_T_1 = gen_small_0_cnt_loop_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_small_0_cnt_loop_ccnt_T_2 = nxt_7 ? 10'h0 : _gen_small_0_cnt_loop_ccnt_T_1; // @[utils.scala 18:20]
  wire  nxt_8 = gen_small_0_cnt_y_ccnt == gen_small_0_cnt_y_cend; // @[utils.scala 17:20]
  wire [9:0] _gen_small_0_cnt_y_ccnt_T_1 = gen_small_0_cnt_y_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_small_0_cnt_y_ccnt_T_2 = nxt_8 ? 10'h0 : _gen_small_0_cnt_y_ccnt_T_1; // @[utils.scala 18:20]
  wire  nxt_9 = ~gen_small_0_cnt_ups_ccnt; // @[utils.scala 17:20]
  wire  _gen_small_0_cnt_ups_ccnt_T_2 = nxt_9 ? 1'h0 : gen_small_0_cnt_ups_ccnt + 1'h1; // @[utils.scala 18:20]
  wire  nxt_10 = gen_small_0_cnt_swap_ccnt == gen_small_0_cnt_swap_cend; // @[utils.scala 17:20]
  wire  _gen_small_0_cnt_swap_ccnt_T_2 = nxt_10 ? 1'h0 : gen_small_0_cnt_swap_ccnt + 1'h1; // @[utils.scala 18:20]
  wire [9:0] _nxt_addr_T_7 = gen_small_0_now_addr + 10'h1; // @[gen_addr.scala 172:53]
  wire [9:0] _GEN_30 = nxt_10 ? _nxt_addr_T_7 : gen_small_0_y_begin_addr; // @[gen_addr.scala 171:49 gen_addr.scala 172:42 gen_addr.scala 175:42]
  wire [9:0] _GEN_33 = nxt_9 ? _GEN_30 : gen_small_0_y_begin_addr; // @[gen_addr.scala 170:44 gen_addr.scala 180:38]
  wire [9:0] _GEN_39 = nxt_8 ? _GEN_33 : _nxt_addr_T_7; // @[gen_addr.scala 169:38 gen_addr.scala 183:34]
  wire [9:0] _GEN_47 = nxt_7 ? _GEN_39 : gen_small_0_ic_begin_addr; // @[gen_addr.scala 168:37 gen_addr.scala 187:30]
  wire [9:0] _GEN_56 = nxt_6 ? _GEN_47 : _nxt_addr_T_7; // @[gen_addr.scala 167:31 gen_addr.scala 190:26]
  wire [9:0] nxt_addr_1 = nxt_5 | gen_small_0_start ? _GEN_56 : 10'h0; // @[gen_addr.scala 165:39 gen_addr.scala 164:18]
  wire [9:0] _gen_small_0_y_begin_addr_nxt_T_1 = nxt_addr_1 - gen_small_0_max_addr; // @[gen_addr.scala 49:24]
  wire [10:0] _gen_small_0_y_begin_addr_nxt_T_2 = {{1'd0}, _gen_small_0_y_begin_addr_nxt_T_1}; // @[gen_addr.scala 49:33]
  wire [9:0] gen_small_0_y_begin_addr_nxt = nxt_addr_1 >= gen_small_0_max_addr ? _gen_small_0_y_begin_addr_nxt_T_2[9:0]
     : nxt_addr_1; // @[gen_addr.scala 48:29 gen_addr.scala 49:17 gen_addr.scala 51:17]
  wire [9:0] _GEN_31 = nxt_10 ? gen_small_0_y_begin_addr_nxt : gen_small_0_y_begin_addr; // @[gen_addr.scala 171:49 gen_addr.scala 173:46 read.scala 26:22]
  wire  _GEN_32 = nxt_9 ? _gen_small_0_cnt_swap_ccnt_T_2 : gen_small_0_cnt_swap_ccnt; // @[gen_addr.scala 170:44 utils.scala 18:14 read.scala 26:22]
  wire [9:0] _GEN_34 = nxt_9 ? _GEN_31 : gen_small_0_y_begin_addr; // @[gen_addr.scala 170:44 read.scala 26:22]
  wire  _GEN_37 = nxt_8 ? _gen_small_0_cnt_ups_ccnt_T_2 : gen_small_0_cnt_ups_ccnt; // @[gen_addr.scala 169:38 utils.scala 18:14 read.scala 26:22]
  wire  _GEN_38 = nxt_8 ? _GEN_32 : gen_small_0_cnt_swap_ccnt; // @[gen_addr.scala 169:38 read.scala 26:22]
  wire [9:0] _GEN_40 = nxt_8 ? _GEN_34 : gen_small_0_y_begin_addr; // @[gen_addr.scala 169:38 read.scala 26:22]
  wire [9:0] _GEN_44 = nxt_7 ? _gen_small_0_cnt_y_ccnt_T_2 : gen_small_0_cnt_y_ccnt; // @[gen_addr.scala 168:37 utils.scala 18:14 read.scala 26:22]
  wire  _GEN_45 = nxt_7 ? _GEN_37 : gen_small_0_cnt_ups_ccnt; // @[gen_addr.scala 168:37 read.scala 26:22]
  wire  _GEN_46 = nxt_7 ? _GEN_38 : gen_small_0_cnt_swap_ccnt; // @[gen_addr.scala 168:37 read.scala 26:22]
  wire [9:0] _GEN_48 = nxt_7 ? _GEN_40 : gen_small_0_y_begin_addr; // @[gen_addr.scala 168:37 read.scala 26:22]
  wire [9:0] _GEN_51 = nxt_7 ? gen_small_0_y_begin_addr_nxt : gen_small_0_ic_begin_addr; // @[gen_addr.scala 168:37 gen_addr.scala 185:35 read.scala 26:22]
  wire [9:0] _GEN_52 = nxt_6 ? _gen_small_0_cnt_loop_ccnt_T_2 : gen_small_0_cnt_loop_ccnt; // @[gen_addr.scala 167:31 utils.scala 18:14 read.scala 26:22]
  wire [9:0] _GEN_53 = nxt_6 ? _GEN_44 : gen_small_0_cnt_y_ccnt; // @[gen_addr.scala 167:31 read.scala 26:22]
  wire  _GEN_54 = nxt_6 ? _GEN_45 : gen_small_0_cnt_ups_ccnt; // @[gen_addr.scala 167:31 read.scala 26:22]
  wire  _GEN_55 = nxt_6 ? _GEN_46 : gen_small_0_cnt_swap_ccnt; // @[gen_addr.scala 167:31 read.scala 26:22]
  wire [9:0] _GEN_57 = nxt_6 ? _GEN_48 : gen_small_0_y_begin_addr; // @[gen_addr.scala 167:31 read.scala 26:22]
  wire [9:0] _GEN_60 = nxt_6 ? _GEN_51 : gen_small_0_ic_begin_addr; // @[gen_addr.scala 167:31 read.scala 26:22]
  wire  _GEN_62 = nxt_5 | gen_small_0_start | gen_small_0_start; // @[gen_addr.scala 165:39 gen_addr.scala 166:19 read.scala 26:22]
  wire  _GEN_402 = io_valid_in & ~gen_big_flag_end; // @[read.scala 31:28 read.scala 40:22 read.scala 21:18]
  wire [2:0] _GEN_403 = io_valid_in ? gen_big_bank_id : 3'h0; // @[read.scala 31:28 read.scala 41:21 read.scala 22:17]
  wire [9:0] _GEN_406 = io_valid_in ? gen_small_0_now_addr : 10'h0; // @[read.scala 31:28 read.scala 41:21 read.scala 22:17]
  wire  _GEN_454 = io_flag_job | gen_small_0_cnt_swap_cend; // @[read.scala 28:22 utils.scala 22:14 read.scala 26:22]
  assign io_valid_out = io_flag_job ? 1'h0 : _GEN_402; // @[read.scala 28:22 read.scala 21:18]
  assign io_to_banks_addrs_0_bank_id = io_flag_job ? 3'h0 : _GEN_403; // @[read.scala 28:22 read.scala 22:17]
  assign io_to_banks_addrs_1_addr = io_flag_job ? 10'h0 : _GEN_406; // @[read.scala 28:22 read.scala 22:17]
  always @(posedge clock) begin
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_ic_ccnt <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt) begin // @[utils.scala 18:20]
        gen_big_cnt_ic_ccnt <= 10'h0;
      end else begin
        gen_big_cnt_ic_ccnt <= _gen_big_cnt_ic_ccnt_T_1;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_ic_cend <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_ic_cend <= io_job_big_cnt_ic_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_x_ccnt <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_x_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt) begin // @[gen_addr.scala 81:27]
        gen_big_cnt_x_ccnt <= _GEN_15;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_x_cend <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_x_cend <= io_job_big_cnt_x_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_y_ccnt <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_y_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt) begin // @[gen_addr.scala 81:27]
        gen_big_cnt_y_ccnt <= _GEN_13;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_y_cend <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_y_cend <= io_job_big_cnt_y_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_bank_id <= 3'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_bank_id <= io_job_big_bank_id; // @[gen_addr.scala 64:17]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_loop_ccnt <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_loop_ccnt <= io_job_big_begin_loop; // @[utils.scala 27:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt) begin // @[gen_addr.scala 81:27]
        gen_big_cnt_loop_ccnt <= _gen_big_cnt_loop_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_loop_cend <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_loop_cend <= io_job_big_cnt_loop_end; // @[utils.scala 26:14]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_cnt_ups_ccnt <= 1'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_big_cnt_ups_ccnt <= 1'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt) begin // @[gen_addr.scala 81:27]
        gen_big_cnt_ups_ccnt <= _GEN_14;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_big_flag_end <= 1'h0; // @[read.scala 26:22]
    end else if (!(io_flag_job)) begin // @[read.scala 28:22]
      if (io_valid_in) begin // @[read.scala 31:28]
        if (nxt) begin // @[gen_addr.scala 81:27]
          gen_big_flag_end <= _GEN_16;
        end
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_max_addr <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_max_addr <= io_job_small_0_max_addr; // @[gen_addr.scala 56:18]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_now_addr <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_now_addr <= 10'h0; // @[gen_addr.scala 58:18]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5 | gen_small_0_start) begin // @[gen_addr.scala 165:39]
        gen_small_0_now_addr <= gen_small_0_y_begin_addr_nxt; // @[gen_addr.scala 192:22]
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_ic_ccnt <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5 | gen_small_0_start) begin // @[gen_addr.scala 165:39]
        gen_small_0_cnt_ic_ccnt <= _gen_small_0_cnt_ic_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_ic_cend <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_ic_cend <= io_job_small_0_cnt_ic_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_y_ccnt <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_y_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5 | gen_small_0_start) begin // @[gen_addr.scala 165:39]
        gen_small_0_cnt_y_ccnt <= _GEN_53;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_y_cend <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_y_cend <= io_job_small_0_cnt_y_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_invalid_ccnt <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_invalid_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5) begin // @[utils.scala 18:20]
        gen_small_0_cnt_invalid_ccnt <= 10'h0;
      end else begin
        gen_small_0_cnt_invalid_ccnt <= _gen_small_0_cnt_invalid_ccnt_T_1;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_invalid_cend <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_invalid_cend <= io_job_small_0_cnt_invalid_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_ups_ccnt <= 1'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_ups_ccnt <= 1'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5 | gen_small_0_start) begin // @[gen_addr.scala 165:39]
        gen_small_0_cnt_ups_ccnt <= _GEN_54;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_loop_ccnt <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_loop_ccnt <= io_job_small_0_begin_loop; // @[utils.scala 27:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5 | gen_small_0_start) begin // @[gen_addr.scala 165:39]
        gen_small_0_cnt_loop_ccnt <= _GEN_52;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_loop_cend <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_loop_cend <= io_job_small_0_cnt_loop_end; // @[utils.scala 26:14]
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_swap_ccnt <= 1'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_cnt_swap_ccnt <= 1'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5 | gen_small_0_start) begin // @[gen_addr.scala 165:39]
        gen_small_0_cnt_swap_ccnt <= _GEN_55;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_cnt_swap_cend <= 1'h0; // @[read.scala 26:22]
    end else begin
      gen_small_0_cnt_swap_cend <= _GEN_454;
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_y_begin_addr <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_y_begin_addr <= 10'h0; // @[gen_addr.scala 235:22]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5 | gen_small_0_start) begin // @[gen_addr.scala 165:39]
        gen_small_0_y_begin_addr <= _GEN_57;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_ic_begin_addr <= 10'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_ic_begin_addr <= 10'h0; // @[gen_addr.scala 236:23]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      if (nxt_5 | gen_small_0_start) begin // @[gen_addr.scala 165:39]
        gen_small_0_ic_begin_addr <= _GEN_60;
      end
    end
    if (reset) begin // @[read.scala 26:22]
      gen_small_0_start <= 1'h0; // @[read.scala 26:22]
    end else if (io_flag_job) begin // @[read.scala 28:22]
      gen_small_0_start <= 1'h0; // @[gen_addr.scala 234:15]
    end else if (io_valid_in) begin // @[read.scala 31:28]
      gen_small_0_start <= _GEN_62;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  gen_big_cnt_ic_ccnt = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  gen_big_cnt_ic_cend = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  gen_big_cnt_x_ccnt = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  gen_big_cnt_x_cend = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  gen_big_cnt_y_ccnt = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  gen_big_cnt_y_cend = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  gen_big_bank_id = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  gen_big_cnt_loop_ccnt = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  gen_big_cnt_loop_cend = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  gen_big_cnt_ups_ccnt = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  gen_big_flag_end = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  gen_small_0_max_addr = _RAND_11[9:0];
  _RAND_12 = {1{`RANDOM}};
  gen_small_0_now_addr = _RAND_12[9:0];
  _RAND_13 = {1{`RANDOM}};
  gen_small_0_cnt_ic_ccnt = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  gen_small_0_cnt_ic_cend = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  gen_small_0_cnt_y_ccnt = _RAND_15[9:0];
  _RAND_16 = {1{`RANDOM}};
  gen_small_0_cnt_y_cend = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  gen_small_0_cnt_invalid_ccnt = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  gen_small_0_cnt_invalid_cend = _RAND_18[9:0];
  _RAND_19 = {1{`RANDOM}};
  gen_small_0_cnt_ups_ccnt = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  gen_small_0_cnt_loop_ccnt = _RAND_20[9:0];
  _RAND_21 = {1{`RANDOM}};
  gen_small_0_cnt_loop_cend = _RAND_21[9:0];
  _RAND_22 = {1{`RANDOM}};
  gen_small_0_cnt_swap_ccnt = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  gen_small_0_cnt_swap_cend = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  gen_small_0_y_begin_addr = _RAND_24[9:0];
  _RAND_25 = {1{`RANDOM}};
  gen_small_0_ic_begin_addr = _RAND_25[9:0];
  _RAND_26 = {1{`RANDOM}};
  gen_small_0_start = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PackReadData(
  input         clock,
  input         reset,
  input         io_valid_in,
  output        io_valid_out,
  input         io_flag_job,
  input  [9:0]  io_job_cnt_x_end,
  input  [9:0]  io_job_cnt_y_end,
  input  [9:0]  io_job_in_chan,
  input  [15:0] io_from_big_0_data_0,
  input  [15:0] io_from_big_0_data_1,
  input  [15:0] io_from_big_0_data_2,
  input  [15:0] io_from_big_0_data_3,
  input  [15:0] io_from_big_0_data_4,
  input  [15:0] io_from_big_0_data_5,
  input  [15:0] io_from_big_0_data_6,
  input  [15:0] io_from_big_0_data_7,
  input  [15:0] io_from_big_0_data_8,
  input  [15:0] io_from_big_0_data_9,
  input  [15:0] io_from_big_0_data_10,
  input  [15:0] io_from_big_0_data_11,
  input  [15:0] io_from_big_0_data_12,
  input  [15:0] io_from_big_0_data_13,
  input  [15:0] io_from_big_0_data_14,
  input  [15:0] io_from_big_0_data_15,
  input  [15:0] io_from_big_0_data_16,
  input  [15:0] io_from_big_0_data_17,
  input  [15:0] io_from_big_0_data_18,
  input  [15:0] io_from_big_0_data_19,
  input  [15:0] io_from_big_0_data_20,
  input  [15:0] io_from_big_0_data_21,
  input  [15:0] io_from_big_0_data_22,
  input  [15:0] io_from_big_0_data_23,
  input  [15:0] io_from_big_0_data_24,
  input  [15:0] io_from_big_0_data_25,
  input  [15:0] io_from_big_0_data_26,
  input  [15:0] io_from_big_0_data_27,
  input  [15:0] io_from_big_0_data_28,
  input  [15:0] io_from_big_0_data_29,
  input  [15:0] io_from_big_0_data_30,
  input  [15:0] io_from_big_0_data_31,
  input  [15:0] io_from_big_0_data_32,
  input  [15:0] io_from_big_0_data_33,
  input  [15:0] io_from_big_0_data_34,
  input  [15:0] io_from_big_0_data_35,
  input  [15:0] io_from_big_0_data_36,
  input  [15:0] io_from_big_0_data_37,
  input  [15:0] io_from_big_0_data_38,
  input  [15:0] io_from_big_0_data_39,
  input  [15:0] io_from_big_0_data_40,
  input  [15:0] io_from_big_0_data_41,
  input  [15:0] io_from_big_0_data_42,
  input  [15:0] io_from_big_0_data_43,
  input  [15:0] io_from_big_0_data_44,
  input  [15:0] io_from_big_0_data_45,
  input  [15:0] io_from_big_0_data_46,
  input  [15:0] io_from_big_0_data_47,
  input  [15:0] io_from_big_1_data_0,
  input  [15:0] io_from_big_1_data_1,
  input  [15:0] io_from_big_1_data_2,
  input  [15:0] io_from_big_1_data_3,
  input  [15:0] io_from_big_1_data_4,
  input  [15:0] io_from_big_1_data_5,
  input  [15:0] io_from_big_1_data_6,
  input  [15:0] io_from_big_1_data_7,
  input  [15:0] io_from_big_1_data_8,
  input  [15:0] io_from_big_1_data_9,
  input  [15:0] io_from_big_1_data_10,
  input  [15:0] io_from_big_1_data_11,
  input  [15:0] io_from_big_1_data_12,
  input  [15:0] io_from_big_1_data_13,
  input  [15:0] io_from_big_1_data_14,
  input  [15:0] io_from_big_1_data_15,
  input  [15:0] io_from_big_1_data_16,
  input  [15:0] io_from_big_1_data_17,
  input  [15:0] io_from_big_1_data_18,
  input  [15:0] io_from_big_1_data_19,
  input  [15:0] io_from_big_1_data_20,
  input  [15:0] io_from_big_1_data_21,
  input  [15:0] io_from_big_1_data_22,
  input  [15:0] io_from_big_1_data_23,
  input  [15:0] io_from_big_1_data_24,
  input  [15:0] io_from_big_1_data_25,
  input  [15:0] io_from_big_1_data_26,
  input  [15:0] io_from_big_1_data_27,
  input  [15:0] io_from_big_1_data_28,
  input  [15:0] io_from_big_1_data_29,
  input  [15:0] io_from_big_1_data_30,
  input  [15:0] io_from_big_1_data_31,
  input  [15:0] io_from_big_1_data_32,
  input  [15:0] io_from_big_1_data_33,
  input  [15:0] io_from_big_1_data_34,
  input  [15:0] io_from_big_1_data_35,
  input  [15:0] io_from_big_1_data_36,
  input  [15:0] io_from_big_1_data_37,
  input  [15:0] io_from_big_1_data_38,
  input  [15:0] io_from_big_1_data_39,
  input  [15:0] io_from_big_1_data_40,
  input  [15:0] io_from_big_1_data_41,
  input  [15:0] io_from_big_1_data_42,
  input  [15:0] io_from_big_1_data_43,
  input  [15:0] io_from_big_1_data_44,
  input  [15:0] io_from_big_1_data_45,
  input  [15:0] io_from_big_1_data_46,
  input  [15:0] io_from_big_1_data_47,
  input  [15:0] io_from_small_0_0_data_0,
  input  [15:0] io_from_small_0_0_data_1,
  input  [15:0] io_from_small_0_0_data_2,
  input  [15:0] io_from_small_0_0_data_3,
  input  [15:0] io_from_small_0_0_data_4,
  input  [15:0] io_from_small_0_0_data_5,
  input  [15:0] io_from_small_0_0_data_6,
  input  [15:0] io_from_small_0_0_data_7,
  input  [15:0] io_from_small_0_1_data_0,
  input  [15:0] io_from_small_0_1_data_1,
  input  [15:0] io_from_small_0_1_data_2,
  input  [15:0] io_from_small_0_1_data_3,
  input  [15:0] io_from_small_0_1_data_4,
  input  [15:0] io_from_small_0_1_data_5,
  input  [15:0] io_from_small_0_1_data_6,
  input  [15:0] io_from_small_0_1_data_7,
  input  [15:0] io_from_small_0_2_data_0,
  input  [15:0] io_from_small_0_2_data_1,
  input  [15:0] io_from_small_0_2_data_2,
  input  [15:0] io_from_small_0_2_data_3,
  input  [15:0] io_from_small_0_2_data_4,
  input  [15:0] io_from_small_0_2_data_5,
  input  [15:0] io_from_small_0_2_data_6,
  input  [15:0] io_from_small_0_2_data_7,
  input  [15:0] io_from_small_0_3_data_0,
  input  [15:0] io_from_small_0_3_data_1,
  input  [15:0] io_from_small_0_3_data_2,
  input  [15:0] io_from_small_0_3_data_3,
  input  [15:0] io_from_small_0_3_data_4,
  input  [15:0] io_from_small_0_3_data_5,
  input  [15:0] io_from_small_0_3_data_6,
  input  [15:0] io_from_small_0_3_data_7,
  input  [15:0] io_from_small_1_0_data_0,
  input  [15:0] io_from_small_1_0_data_1,
  input  [15:0] io_from_small_1_0_data_2,
  input  [15:0] io_from_small_1_0_data_3,
  input  [15:0] io_from_small_1_0_data_4,
  input  [15:0] io_from_small_1_0_data_5,
  input  [15:0] io_from_small_1_0_data_6,
  input  [15:0] io_from_small_1_0_data_7,
  input  [15:0] io_from_small_1_1_data_0,
  input  [15:0] io_from_small_1_1_data_1,
  input  [15:0] io_from_small_1_1_data_2,
  input  [15:0] io_from_small_1_1_data_3,
  input  [15:0] io_from_small_1_1_data_4,
  input  [15:0] io_from_small_1_1_data_5,
  input  [15:0] io_from_small_1_1_data_6,
  input  [15:0] io_from_small_1_1_data_7,
  input  [15:0] io_from_small_1_2_data_0,
  input  [15:0] io_from_small_1_2_data_1,
  input  [15:0] io_from_small_1_2_data_2,
  input  [15:0] io_from_small_1_2_data_3,
  input  [15:0] io_from_small_1_2_data_4,
  input  [15:0] io_from_small_1_2_data_5,
  input  [15:0] io_from_small_1_2_data_6,
  input  [15:0] io_from_small_1_2_data_7,
  input  [15:0] io_from_small_1_3_data_0,
  input  [15:0] io_from_small_1_3_data_1,
  input  [15:0] io_from_small_1_3_data_2,
  input  [15:0] io_from_small_1_3_data_3,
  input  [15:0] io_from_small_1_3_data_4,
  input  [15:0] io_from_small_1_3_data_5,
  input  [15:0] io_from_small_1_3_data_6,
  input  [15:0] io_from_small_1_3_data_7,
  output [15:0] io_output_mat_0,
  output [15:0] io_output_mat_1,
  output [15:0] io_output_mat_2,
  output [15:0] io_output_mat_3,
  output [15:0] io_output_mat_4,
  output [15:0] io_output_mat_5,
  output [15:0] io_output_mat_6,
  output [15:0] io_output_mat_7,
  output [15:0] io_output_mat_8,
  output [15:0] io_output_mat_9,
  output [15:0] io_output_mat_10,
  output [15:0] io_output_mat_11,
  output [15:0] io_output_mat_12,
  output [15:0] io_output_mat_13,
  output [15:0] io_output_mat_14,
  output [15:0] io_output_mat_15,
  output [15:0] io_output_mat_16,
  output [15:0] io_output_mat_17,
  output [15:0] io_output_mat_18,
  output [15:0] io_output_mat_19,
  output [15:0] io_output_mat_20,
  output [15:0] io_output_mat_21,
  output [15:0] io_output_mat_22,
  output [15:0] io_output_mat_23,
  output [15:0] io_output_mat_24,
  output [15:0] io_output_mat_25,
  output [15:0] io_output_mat_26,
  output [15:0] io_output_mat_27,
  output [15:0] io_output_mat_28,
  output [15:0] io_output_mat_29,
  output [15:0] io_output_mat_30,
  output [15:0] io_output_mat_31,
  output [15:0] io_output_mat_32,
  output [15:0] io_output_mat_33,
  output [15:0] io_output_mat_34,
  output [15:0] io_output_mat_35,
  output [15:0] io_output_mat_36,
  output [15:0] io_output_mat_37,
  output [15:0] io_output_mat_38,
  output [15:0] io_output_mat_39,
  output [15:0] io_output_mat_40,
  output [15:0] io_output_mat_41,
  output [15:0] io_output_mat_42,
  output [15:0] io_output_mat_43,
  output [15:0] io_output_mat_44,
  output [15:0] io_output_mat_45,
  output [15:0] io_output_mat_46,
  output [15:0] io_output_mat_47,
  output [15:0] io_output_mat_48,
  output [15:0] io_output_mat_49,
  output [15:0] io_output_mat_50,
  output [15:0] io_output_mat_51,
  output [15:0] io_output_mat_52,
  output [15:0] io_output_mat_53,
  output [15:0] io_output_mat_54,
  output [15:0] io_output_mat_55,
  output [15:0] io_output_mat_56,
  output [15:0] io_output_mat_57,
  output [15:0] io_output_mat_58,
  output [15:0] io_output_mat_59,
  output [15:0] io_output_mat_60,
  output [15:0] io_output_mat_61,
  output [15:0] io_output_mat_62,
  output [15:0] io_output_mat_63,
  output [15:0] io_output_up_0,
  output [15:0] io_output_up_1,
  output [15:0] io_output_up_2,
  output [15:0] io_output_up_3,
  output [15:0] io_output_up_4,
  output [15:0] io_output_up_5,
  output [15:0] io_output_up_6,
  output [15:0] io_output_up_7,
  output [15:0] io_output_up_8,
  output [15:0] io_output_up_9,
  output [15:0] io_output_down_0,
  output [15:0] io_output_down_1,
  output [15:0] io_output_down_2,
  output [15:0] io_output_down_3,
  output [15:0] io_output_down_4,
  output [15:0] io_output_down_5,
  output [15:0] io_output_down_6,
  output [15:0] io_output_down_7,
  output [15:0] io_output_down_8,
  output [15:0] io_output_down_9,
  output [15:0] io_output_left_0,
  output [15:0] io_output_left_1,
  output [15:0] io_output_left_2,
  output [15:0] io_output_left_3,
  output [15:0] io_output_left_4,
  output [15:0] io_output_left_5,
  output [15:0] io_output_left_6,
  output [15:0] io_output_left_7,
  output [15:0] io_output_right_0,
  output [15:0] io_output_right_1,
  output [15:0] io_output_right_2,
  output [15:0] io_output_right_3,
  output [15:0] io_output_right_4,
  output [15:0] io_output_right_5,
  output [15:0] io_output_right_6,
  output [15:0] io_output_right_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] cache_0_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_0_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_1_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_2_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_3_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_4_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_5_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_6_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_7_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_8_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_9_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_10_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_11_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_12_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_13_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_14_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_15_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_16_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_17_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_18_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_19_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_20_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_21_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_22_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_23_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_24_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_25_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_26_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_27_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_28_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_29_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_30_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_31_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_32_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_33_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_34_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_35_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_36_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_37_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_38_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_39_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_40_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_41_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_42_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_43_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_44_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_45_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_46_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_47_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_48_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_49_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_50_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_51_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_52_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_53_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_54_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_55_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_56_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_57_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_58_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_59_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_60_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_61_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_62_9; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_0; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_1; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_2; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_3; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_4; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_5; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_6; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_7; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_8; // @[read_pack.scala 23:24]
  reg [15:0] cache_63_9; // @[read_pack.scala 23:24]
  reg [9:0] cnt_ic_ccnt; // @[read_pack.scala 25:25]
  reg [9:0] cnt_ic_cend; // @[read_pack.scala 25:25]
  reg [9:0] cnt_x_ccnt; // @[read_pack.scala 26:24]
  reg [9:0] cnt_x_cend; // @[read_pack.scala 26:24]
  reg [9:0] cnt_y_ccnt; // @[read_pack.scala 27:24]
  reg [9:0] cnt_y_cend; // @[read_pack.scala 27:24]
  reg  state; // @[read_pack.scala 33:24]
  wire  nxt = cnt_ic_ccnt == cnt_ic_cend; // @[utils.scala 17:20]
  wire [9:0] _cnt_ic_ccnt_T_1 = cnt_ic_ccnt + 10'h1; // @[utils.scala 18:35]
  wire  _state_T = ~state; // @[read_pack.scala 51:22]
  wire  nxt_1 = cnt_y_ccnt == cnt_y_cend; // @[utils.scala 17:20]
  wire [9:0] _cnt_y_ccnt_T_1 = cnt_y_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _cnt_y_ccnt_T_2 = nxt_1 ? 10'h0 : _cnt_y_ccnt_T_1; // @[utils.scala 18:20]
  wire  nxt_2 = cnt_x_ccnt == cnt_x_cend; // @[utils.scala 17:20]
  wire [9:0] _cnt_x_ccnt_T_1 = cnt_x_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _cnt_x_ccnt_T_2 = nxt_2 ? 10'h0 : _cnt_x_ccnt_T_1; // @[utils.scala 18:20]
  wire [9:0] _GEN_0 = nxt_1 ? _cnt_x_ccnt_T_2 : cnt_x_ccnt; // @[read_pack.scala 52:30 utils.scala 18:14 read_pack.scala 26:24]
  wire [15:0] _GEN_5 = state ? $signed(io_from_big_1_data_0) : $signed(io_from_big_0_data_0); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_7 = state ? $signed(io_from_big_1_data_1) : $signed(io_from_big_0_data_1); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_9 = state ? $signed(io_from_big_1_data_2) : $signed(io_from_big_0_data_2); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_11 = state ? $signed(io_from_big_1_data_3) : $signed(io_from_big_0_data_3); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_13 = state ? $signed(io_from_big_1_data_4) : $signed(io_from_big_0_data_4); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_15 = state ? $signed(io_from_big_1_data_5) : $signed(io_from_big_0_data_5); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_17 = state ? $signed(io_from_small_1_1_data_0) : $signed(io_from_small_0_1_data_0); // @[read_pack.scala 39:34 read_pack.scala 39:34]
  wire [15:0] _GEN_19 = state ? $signed(io_from_small_1_2_data_0) : $signed(io_from_small_0_2_data_0); // @[read_pack.scala 40:34 read_pack.scala 40:34]
  wire [15:0] _GEN_21 = state ? $signed(io_from_big_1_data_6) : $signed(io_from_big_0_data_6); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_23 = state ? $signed(io_from_big_1_data_7) : $signed(io_from_big_0_data_7); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_25 = state ? $signed(io_from_big_1_data_8) : $signed(io_from_big_0_data_8); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_27 = state ? $signed(io_from_big_1_data_9) : $signed(io_from_big_0_data_9); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_29 = state ? $signed(io_from_big_1_data_10) : $signed(io_from_big_0_data_10); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_31 = state ? $signed(io_from_big_1_data_11) : $signed(io_from_big_0_data_11); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_33 = state ? $signed(io_from_small_1_1_data_1) : $signed(io_from_small_0_1_data_1); // @[read_pack.scala 39:34 read_pack.scala 39:34]
  wire [15:0] _GEN_35 = state ? $signed(io_from_small_1_2_data_1) : $signed(io_from_small_0_2_data_1); // @[read_pack.scala 40:34 read_pack.scala 40:34]
  wire [15:0] _GEN_37 = state ? $signed(io_from_big_1_data_12) : $signed(io_from_big_0_data_12); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_39 = state ? $signed(io_from_big_1_data_13) : $signed(io_from_big_0_data_13); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_41 = state ? $signed(io_from_big_1_data_14) : $signed(io_from_big_0_data_14); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_43 = state ? $signed(io_from_big_1_data_15) : $signed(io_from_big_0_data_15); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_45 = state ? $signed(io_from_big_1_data_16) : $signed(io_from_big_0_data_16); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_47 = state ? $signed(io_from_big_1_data_17) : $signed(io_from_big_0_data_17); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_49 = state ? $signed(io_from_small_1_1_data_2) : $signed(io_from_small_0_1_data_2); // @[read_pack.scala 39:34 read_pack.scala 39:34]
  wire [15:0] _GEN_51 = state ? $signed(io_from_small_1_2_data_2) : $signed(io_from_small_0_2_data_2); // @[read_pack.scala 40:34 read_pack.scala 40:34]
  wire [15:0] _GEN_53 = state ? $signed(io_from_big_1_data_18) : $signed(io_from_big_0_data_18); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_55 = state ? $signed(io_from_big_1_data_19) : $signed(io_from_big_0_data_19); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_57 = state ? $signed(io_from_big_1_data_20) : $signed(io_from_big_0_data_20); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_59 = state ? $signed(io_from_big_1_data_21) : $signed(io_from_big_0_data_21); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_61 = state ? $signed(io_from_big_1_data_22) : $signed(io_from_big_0_data_22); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_63 = state ? $signed(io_from_big_1_data_23) : $signed(io_from_big_0_data_23); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_65 = state ? $signed(io_from_small_1_1_data_3) : $signed(io_from_small_0_1_data_3); // @[read_pack.scala 39:34 read_pack.scala 39:34]
  wire [15:0] _GEN_67 = state ? $signed(io_from_small_1_2_data_3) : $signed(io_from_small_0_2_data_3); // @[read_pack.scala 40:34 read_pack.scala 40:34]
  wire [15:0] _GEN_69 = state ? $signed(io_from_big_1_data_24) : $signed(io_from_big_0_data_24); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_71 = state ? $signed(io_from_big_1_data_25) : $signed(io_from_big_0_data_25); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_73 = state ? $signed(io_from_big_1_data_26) : $signed(io_from_big_0_data_26); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_75 = state ? $signed(io_from_big_1_data_27) : $signed(io_from_big_0_data_27); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_77 = state ? $signed(io_from_big_1_data_28) : $signed(io_from_big_0_data_28); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_79 = state ? $signed(io_from_big_1_data_29) : $signed(io_from_big_0_data_29); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_81 = state ? $signed(io_from_small_1_1_data_4) : $signed(io_from_small_0_1_data_4); // @[read_pack.scala 39:34 read_pack.scala 39:34]
  wire [15:0] _GEN_83 = state ? $signed(io_from_small_1_2_data_4) : $signed(io_from_small_0_2_data_4); // @[read_pack.scala 40:34 read_pack.scala 40:34]
  wire [15:0] _GEN_85 = state ? $signed(io_from_big_1_data_30) : $signed(io_from_big_0_data_30); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_87 = state ? $signed(io_from_big_1_data_31) : $signed(io_from_big_0_data_31); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_89 = state ? $signed(io_from_big_1_data_32) : $signed(io_from_big_0_data_32); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_91 = state ? $signed(io_from_big_1_data_33) : $signed(io_from_big_0_data_33); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_93 = state ? $signed(io_from_big_1_data_34) : $signed(io_from_big_0_data_34); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_95 = state ? $signed(io_from_big_1_data_35) : $signed(io_from_big_0_data_35); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_97 = state ? $signed(io_from_small_1_1_data_5) : $signed(io_from_small_0_1_data_5); // @[read_pack.scala 39:34 read_pack.scala 39:34]
  wire [15:0] _GEN_99 = state ? $signed(io_from_small_1_2_data_5) : $signed(io_from_small_0_2_data_5); // @[read_pack.scala 40:34 read_pack.scala 40:34]
  wire [15:0] _GEN_101 = state ? $signed(io_from_big_1_data_36) : $signed(io_from_big_0_data_36); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_103 = state ? $signed(io_from_big_1_data_37) : $signed(io_from_big_0_data_37); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_105 = state ? $signed(io_from_big_1_data_38) : $signed(io_from_big_0_data_38); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_107 = state ? $signed(io_from_big_1_data_39) : $signed(io_from_big_0_data_39); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_109 = state ? $signed(io_from_big_1_data_40) : $signed(io_from_big_0_data_40); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_111 = state ? $signed(io_from_big_1_data_41) : $signed(io_from_big_0_data_41); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] _GEN_113 = state ? $signed(io_from_small_1_1_data_6) : $signed(io_from_small_0_1_data_6); // @[read_pack.scala 39:34 read_pack.scala 39:34]
  wire [15:0] _GEN_115 = state ? $signed(io_from_small_1_2_data_6) : $signed(io_from_small_0_2_data_6); // @[read_pack.scala 40:34 read_pack.scala 40:34]
  wire [15:0] nxt_up_2 = state ? $signed(io_from_big_1_data_42) : $signed(io_from_big_0_data_42); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] nxt_up_3 = state ? $signed(io_from_big_1_data_43) : $signed(io_from_big_0_data_43); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] nxt_up_4 = state ? $signed(io_from_big_1_data_44) : $signed(io_from_big_0_data_44); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] nxt_up_5 = state ? $signed(io_from_big_1_data_45) : $signed(io_from_big_0_data_45); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] nxt_up_6 = state ? $signed(io_from_big_1_data_46) : $signed(io_from_big_0_data_46); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] nxt_up_7 = state ? $signed(io_from_big_1_data_47) : $signed(io_from_big_0_data_47); // @[read_pack.scala 38:38 read_pack.scala 38:38]
  wire [15:0] nxt_up_1 = state ? $signed(io_from_small_1_1_data_7) : $signed(io_from_small_0_1_data_7); // @[read_pack.scala 39:34 read_pack.scala 39:34]
  wire [15:0] nxt_up_8 = state ? $signed(io_from_small_1_2_data_7) : $signed(io_from_small_0_2_data_7); // @[read_pack.scala 40:34 read_pack.scala 40:34]
  wire  _T_1 = cnt_x_ccnt == 10'h0; // @[read_pack.scala 62:28]
  wire [15:0] _GEN_133 = state ? $signed(io_from_small_1_0_data_1) : $signed(io_from_small_0_0_data_1); // @[read_pack.scala 65:33 read_pack.scala 65:33]
  wire [15:0] _GEN_134 = cnt_x_ccnt == 10'h0 ? $signed(_GEN_21) : $signed(_GEN_133); // @[read_pack.scala 62:35 read_pack.scala 63:33 read_pack.scala 65:33]
  wire [15:0] _GEN_136 = state ? $signed(io_from_small_1_3_data_1) : $signed(io_from_small_0_3_data_1); // @[read_pack.scala 70:33 read_pack.scala 70:33]
  wire [15:0] _GEN_137 = nxt_2 ? $signed(_GEN_31) : $signed(_GEN_136); // @[read_pack.scala 67:42 read_pack.scala 68:33 read_pack.scala 70:33]
  wire [15:0] _GEN_139 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_0) : $signed(cache_0_0); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_140 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_0) : $signed(_GEN_139); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_141 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_0) : $signed(_GEN_140); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_142 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_0) : $signed(_GEN_141); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_143 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_0) : $signed(_GEN_142); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_144 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_0) : $signed(_GEN_143); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_145 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_0) : $signed(_GEN_144); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_146 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_0) : $signed(_GEN_145); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_147 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_0) : $signed(_GEN_146); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_148 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_0) : $signed(_GEN_147); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_149 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_0) : $signed(_GEN_148); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_150 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_0) : $signed(_GEN_149); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_151 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_0) : $signed(_GEN_150); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_152 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_0) : $signed(_GEN_151); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_153 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_0) : $signed(_GEN_152); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_154 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_0) : $signed(_GEN_153); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_155 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_0) : $signed(_GEN_154); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_156 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_0) : $signed(_GEN_155); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_157 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_0) : $signed(_GEN_156); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_158 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_0) : $signed(_GEN_157); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_159 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_0) : $signed(_GEN_158); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_160 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_0) : $signed(_GEN_159); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_161 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_0) : $signed(_GEN_160); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_162 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_0) : $signed(_GEN_161); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_163 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_0) : $signed(_GEN_162); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_164 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_0) : $signed(_GEN_163); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_165 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_0) : $signed(_GEN_164); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_166 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_0) : $signed(_GEN_165); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_167 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_0) : $signed(_GEN_166); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_168 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_0) : $signed(_GEN_167); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_169 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_0) : $signed(_GEN_168); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_170 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_0) : $signed(_GEN_169); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_171 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_0) : $signed(_GEN_170); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_172 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_0) : $signed(_GEN_171); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_173 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_0) : $signed(_GEN_172); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_174 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_0) : $signed(_GEN_173); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_175 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_0) : $signed(_GEN_174); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_176 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_0) : $signed(_GEN_175); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_177 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_0) : $signed(_GEN_176); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_178 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_0) : $signed(_GEN_177); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_179 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_0) : $signed(_GEN_178); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_180 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_0) : $signed(_GEN_179); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_181 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_0) : $signed(_GEN_180); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_182 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_0) : $signed(_GEN_181); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_183 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_0) : $signed(_GEN_182); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_184 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_0) : $signed(_GEN_183); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_185 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_0) : $signed(_GEN_184); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_186 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_0) : $signed(_GEN_185); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_187 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_0) : $signed(_GEN_186); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_188 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_0) : $signed(_GEN_187); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_189 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_0) : $signed(_GEN_188); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_190 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_0) : $signed(_GEN_189); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_191 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_0) : $signed(_GEN_190); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_192 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_0) : $signed(_GEN_191); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_193 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_0) : $signed(_GEN_192); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_194 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_0) : $signed(_GEN_193); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_195 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_0) : $signed(_GEN_194); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_196 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_0) : $signed(_GEN_195); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_197 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_0) : $signed(_GEN_196); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_198 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_0) : $signed(_GEN_197); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_199 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_0) : $signed(_GEN_198); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_200 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_0) : $signed(_GEN_199); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_201 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_0) : $signed(_GEN_200); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_203 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_1) : $signed(cache_0_1); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_204 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_1) : $signed(_GEN_203); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_205 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_1) : $signed(_GEN_204); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_206 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_1) : $signed(_GEN_205); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_207 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_1) : $signed(_GEN_206); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_208 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_1) : $signed(_GEN_207); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_209 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_1) : $signed(_GEN_208); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_210 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_1) : $signed(_GEN_209); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_211 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_1) : $signed(_GEN_210); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_212 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_1) : $signed(_GEN_211); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_213 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_1) : $signed(_GEN_212); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_214 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_1) : $signed(_GEN_213); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_215 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_1) : $signed(_GEN_214); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_216 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_1) : $signed(_GEN_215); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_217 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_1) : $signed(_GEN_216); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_218 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_1) : $signed(_GEN_217); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_219 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_1) : $signed(_GEN_218); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_220 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_1) : $signed(_GEN_219); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_221 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_1) : $signed(_GEN_220); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_222 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_1) : $signed(_GEN_221); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_223 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_1) : $signed(_GEN_222); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_224 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_1) : $signed(_GEN_223); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_225 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_1) : $signed(_GEN_224); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_226 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_1) : $signed(_GEN_225); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_227 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_1) : $signed(_GEN_226); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_228 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_1) : $signed(_GEN_227); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_229 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_1) : $signed(_GEN_228); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_230 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_1) : $signed(_GEN_229); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_231 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_1) : $signed(_GEN_230); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_232 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_1) : $signed(_GEN_231); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_233 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_1) : $signed(_GEN_232); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_234 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_1) : $signed(_GEN_233); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_235 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_1) : $signed(_GEN_234); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_236 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_1) : $signed(_GEN_235); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_237 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_1) : $signed(_GEN_236); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_238 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_1) : $signed(_GEN_237); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_239 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_1) : $signed(_GEN_238); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_240 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_1) : $signed(_GEN_239); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_241 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_1) : $signed(_GEN_240); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_242 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_1) : $signed(_GEN_241); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_243 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_1) : $signed(_GEN_242); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_244 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_1) : $signed(_GEN_243); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_245 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_1) : $signed(_GEN_244); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_246 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_1) : $signed(_GEN_245); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_247 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_1) : $signed(_GEN_246); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_248 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_1) : $signed(_GEN_247); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_249 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_1) : $signed(_GEN_248); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_250 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_1) : $signed(_GEN_249); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_251 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_1) : $signed(_GEN_250); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_252 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_1) : $signed(_GEN_251); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_253 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_1) : $signed(_GEN_252); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_254 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_1) : $signed(_GEN_253); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_255 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_1) : $signed(_GEN_254); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_256 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_1) : $signed(_GEN_255); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_257 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_1) : $signed(_GEN_256); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_258 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_1) : $signed(_GEN_257); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_259 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_1) : $signed(_GEN_258); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_260 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_1) : $signed(_GEN_259); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_261 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_1) : $signed(_GEN_260); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_262 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_1) : $signed(_GEN_261); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_263 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_1) : $signed(_GEN_262); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_264 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_1) : $signed(_GEN_263); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_265 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_1) : $signed(_GEN_264); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_267 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_2) : $signed(cache_0_2); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_268 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_2) : $signed(_GEN_267); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_269 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_2) : $signed(_GEN_268); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_270 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_2) : $signed(_GEN_269); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_271 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_2) : $signed(_GEN_270); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_272 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_2) : $signed(_GEN_271); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_273 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_2) : $signed(_GEN_272); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_274 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_2) : $signed(_GEN_273); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_275 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_2) : $signed(_GEN_274); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_276 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_2) : $signed(_GEN_275); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_277 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_2) : $signed(_GEN_276); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_278 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_2) : $signed(_GEN_277); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_279 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_2) : $signed(_GEN_278); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_280 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_2) : $signed(_GEN_279); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_281 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_2) : $signed(_GEN_280); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_282 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_2) : $signed(_GEN_281); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_283 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_2) : $signed(_GEN_282); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_284 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_2) : $signed(_GEN_283); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_285 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_2) : $signed(_GEN_284); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_286 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_2) : $signed(_GEN_285); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_287 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_2) : $signed(_GEN_286); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_288 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_2) : $signed(_GEN_287); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_289 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_2) : $signed(_GEN_288); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_290 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_2) : $signed(_GEN_289); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_291 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_2) : $signed(_GEN_290); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_292 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_2) : $signed(_GEN_291); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_293 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_2) : $signed(_GEN_292); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_294 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_2) : $signed(_GEN_293); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_295 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_2) : $signed(_GEN_294); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_296 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_2) : $signed(_GEN_295); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_297 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_2) : $signed(_GEN_296); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_298 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_2) : $signed(_GEN_297); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_299 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_2) : $signed(_GEN_298); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_300 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_2) : $signed(_GEN_299); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_301 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_2) : $signed(_GEN_300); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_302 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_2) : $signed(_GEN_301); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_303 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_2) : $signed(_GEN_302); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_304 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_2) : $signed(_GEN_303); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_305 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_2) : $signed(_GEN_304); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_306 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_2) : $signed(_GEN_305); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_307 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_2) : $signed(_GEN_306); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_308 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_2) : $signed(_GEN_307); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_309 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_2) : $signed(_GEN_308); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_310 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_2) : $signed(_GEN_309); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_311 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_2) : $signed(_GEN_310); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_312 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_2) : $signed(_GEN_311); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_313 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_2) : $signed(_GEN_312); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_314 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_2) : $signed(_GEN_313); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_315 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_2) : $signed(_GEN_314); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_316 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_2) : $signed(_GEN_315); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_317 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_2) : $signed(_GEN_316); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_318 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_2) : $signed(_GEN_317); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_319 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_2) : $signed(_GEN_318); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_320 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_2) : $signed(_GEN_319); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_321 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_2) : $signed(_GEN_320); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_322 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_2) : $signed(_GEN_321); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_323 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_2) : $signed(_GEN_322); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_324 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_2) : $signed(_GEN_323); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_325 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_2) : $signed(_GEN_324); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_326 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_2) : $signed(_GEN_325); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_327 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_2) : $signed(_GEN_326); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_328 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_2) : $signed(_GEN_327); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_329 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_2) : $signed(_GEN_328); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_331 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_3) : $signed(cache_0_3); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_332 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_3) : $signed(_GEN_331); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_333 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_3) : $signed(_GEN_332); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_334 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_3) : $signed(_GEN_333); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_335 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_3) : $signed(_GEN_334); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_336 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_3) : $signed(_GEN_335); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_337 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_3) : $signed(_GEN_336); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_338 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_3) : $signed(_GEN_337); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_339 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_3) : $signed(_GEN_338); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_340 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_3) : $signed(_GEN_339); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_341 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_3) : $signed(_GEN_340); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_342 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_3) : $signed(_GEN_341); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_343 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_3) : $signed(_GEN_342); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_344 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_3) : $signed(_GEN_343); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_345 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_3) : $signed(_GEN_344); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_346 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_3) : $signed(_GEN_345); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_347 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_3) : $signed(_GEN_346); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_348 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_3) : $signed(_GEN_347); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_349 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_3) : $signed(_GEN_348); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_350 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_3) : $signed(_GEN_349); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_351 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_3) : $signed(_GEN_350); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_352 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_3) : $signed(_GEN_351); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_353 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_3) : $signed(_GEN_352); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_354 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_3) : $signed(_GEN_353); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_355 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_3) : $signed(_GEN_354); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_356 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_3) : $signed(_GEN_355); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_357 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_3) : $signed(_GEN_356); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_358 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_3) : $signed(_GEN_357); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_359 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_3) : $signed(_GEN_358); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_360 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_3) : $signed(_GEN_359); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_361 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_3) : $signed(_GEN_360); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_362 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_3) : $signed(_GEN_361); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_363 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_3) : $signed(_GEN_362); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_364 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_3) : $signed(_GEN_363); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_365 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_3) : $signed(_GEN_364); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_366 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_3) : $signed(_GEN_365); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_367 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_3) : $signed(_GEN_366); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_368 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_3) : $signed(_GEN_367); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_369 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_3) : $signed(_GEN_368); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_370 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_3) : $signed(_GEN_369); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_371 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_3) : $signed(_GEN_370); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_372 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_3) : $signed(_GEN_371); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_373 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_3) : $signed(_GEN_372); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_374 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_3) : $signed(_GEN_373); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_375 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_3) : $signed(_GEN_374); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_376 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_3) : $signed(_GEN_375); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_377 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_3) : $signed(_GEN_376); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_378 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_3) : $signed(_GEN_377); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_379 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_3) : $signed(_GEN_378); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_380 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_3) : $signed(_GEN_379); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_381 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_3) : $signed(_GEN_380); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_382 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_3) : $signed(_GEN_381); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_383 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_3) : $signed(_GEN_382); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_384 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_3) : $signed(_GEN_383); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_385 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_3) : $signed(_GEN_384); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_386 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_3) : $signed(_GEN_385); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_387 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_3) : $signed(_GEN_386); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_388 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_3) : $signed(_GEN_387); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_389 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_3) : $signed(_GEN_388); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_390 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_3) : $signed(_GEN_389); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_391 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_3) : $signed(_GEN_390); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_392 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_3) : $signed(_GEN_391); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_393 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_3) : $signed(_GEN_392); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_395 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_4) : $signed(cache_0_4); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_396 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_4) : $signed(_GEN_395); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_397 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_4) : $signed(_GEN_396); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_398 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_4) : $signed(_GEN_397); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_399 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_4) : $signed(_GEN_398); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_400 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_4) : $signed(_GEN_399); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_401 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_4) : $signed(_GEN_400); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_402 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_4) : $signed(_GEN_401); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_403 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_4) : $signed(_GEN_402); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_404 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_4) : $signed(_GEN_403); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_405 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_4) : $signed(_GEN_404); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_406 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_4) : $signed(_GEN_405); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_407 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_4) : $signed(_GEN_406); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_408 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_4) : $signed(_GEN_407); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_409 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_4) : $signed(_GEN_408); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_410 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_4) : $signed(_GEN_409); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_411 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_4) : $signed(_GEN_410); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_412 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_4) : $signed(_GEN_411); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_413 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_4) : $signed(_GEN_412); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_414 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_4) : $signed(_GEN_413); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_415 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_4) : $signed(_GEN_414); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_416 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_4) : $signed(_GEN_415); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_417 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_4) : $signed(_GEN_416); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_418 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_4) : $signed(_GEN_417); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_419 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_4) : $signed(_GEN_418); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_420 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_4) : $signed(_GEN_419); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_421 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_4) : $signed(_GEN_420); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_422 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_4) : $signed(_GEN_421); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_423 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_4) : $signed(_GEN_422); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_424 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_4) : $signed(_GEN_423); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_425 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_4) : $signed(_GEN_424); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_426 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_4) : $signed(_GEN_425); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_427 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_4) : $signed(_GEN_426); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_428 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_4) : $signed(_GEN_427); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_429 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_4) : $signed(_GEN_428); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_430 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_4) : $signed(_GEN_429); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_431 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_4) : $signed(_GEN_430); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_432 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_4) : $signed(_GEN_431); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_433 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_4) : $signed(_GEN_432); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_434 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_4) : $signed(_GEN_433); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_435 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_4) : $signed(_GEN_434); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_436 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_4) : $signed(_GEN_435); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_437 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_4) : $signed(_GEN_436); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_438 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_4) : $signed(_GEN_437); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_439 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_4) : $signed(_GEN_438); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_440 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_4) : $signed(_GEN_439); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_441 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_4) : $signed(_GEN_440); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_442 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_4) : $signed(_GEN_441); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_443 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_4) : $signed(_GEN_442); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_444 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_4) : $signed(_GEN_443); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_445 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_4) : $signed(_GEN_444); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_446 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_4) : $signed(_GEN_445); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_447 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_4) : $signed(_GEN_446); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_448 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_4) : $signed(_GEN_447); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_449 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_4) : $signed(_GEN_448); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_450 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_4) : $signed(_GEN_449); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_451 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_4) : $signed(_GEN_450); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_452 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_4) : $signed(_GEN_451); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_453 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_4) : $signed(_GEN_452); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_454 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_4) : $signed(_GEN_453); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_455 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_4) : $signed(_GEN_454); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_456 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_4) : $signed(_GEN_455); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_457 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_4) : $signed(_GEN_456); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_459 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_5) : $signed(cache_0_5); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_460 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_5) : $signed(_GEN_459); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_461 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_5) : $signed(_GEN_460); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_462 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_5) : $signed(_GEN_461); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_463 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_5) : $signed(_GEN_462); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_464 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_5) : $signed(_GEN_463); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_465 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_5) : $signed(_GEN_464); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_466 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_5) : $signed(_GEN_465); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_467 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_5) : $signed(_GEN_466); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_468 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_5) : $signed(_GEN_467); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_469 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_5) : $signed(_GEN_468); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_470 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_5) : $signed(_GEN_469); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_471 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_5) : $signed(_GEN_470); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_472 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_5) : $signed(_GEN_471); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_473 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_5) : $signed(_GEN_472); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_474 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_5) : $signed(_GEN_473); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_475 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_5) : $signed(_GEN_474); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_476 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_5) : $signed(_GEN_475); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_477 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_5) : $signed(_GEN_476); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_478 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_5) : $signed(_GEN_477); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_479 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_5) : $signed(_GEN_478); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_480 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_5) : $signed(_GEN_479); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_481 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_5) : $signed(_GEN_480); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_482 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_5) : $signed(_GEN_481); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_483 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_5) : $signed(_GEN_482); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_484 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_5) : $signed(_GEN_483); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_485 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_5) : $signed(_GEN_484); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_486 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_5) : $signed(_GEN_485); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_487 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_5) : $signed(_GEN_486); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_488 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_5) : $signed(_GEN_487); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_489 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_5) : $signed(_GEN_488); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_490 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_5) : $signed(_GEN_489); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_491 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_5) : $signed(_GEN_490); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_492 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_5) : $signed(_GEN_491); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_493 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_5) : $signed(_GEN_492); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_494 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_5) : $signed(_GEN_493); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_495 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_5) : $signed(_GEN_494); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_496 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_5) : $signed(_GEN_495); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_497 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_5) : $signed(_GEN_496); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_498 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_5) : $signed(_GEN_497); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_499 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_5) : $signed(_GEN_498); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_500 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_5) : $signed(_GEN_499); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_501 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_5) : $signed(_GEN_500); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_502 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_5) : $signed(_GEN_501); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_503 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_5) : $signed(_GEN_502); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_504 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_5) : $signed(_GEN_503); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_505 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_5) : $signed(_GEN_504); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_506 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_5) : $signed(_GEN_505); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_507 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_5) : $signed(_GEN_506); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_508 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_5) : $signed(_GEN_507); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_509 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_5) : $signed(_GEN_508); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_510 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_5) : $signed(_GEN_509); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_511 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_5) : $signed(_GEN_510); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_512 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_5) : $signed(_GEN_511); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_513 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_5) : $signed(_GEN_512); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_514 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_5) : $signed(_GEN_513); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_515 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_5) : $signed(_GEN_514); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_516 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_5) : $signed(_GEN_515); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_517 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_5) : $signed(_GEN_516); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_518 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_5) : $signed(_GEN_517); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_519 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_5) : $signed(_GEN_518); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_520 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_5) : $signed(_GEN_519); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_521 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_5) : $signed(_GEN_520); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_523 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_6) : $signed(cache_0_6); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_524 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_6) : $signed(_GEN_523); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_525 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_6) : $signed(_GEN_524); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_526 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_6) : $signed(_GEN_525); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_527 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_6) : $signed(_GEN_526); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_528 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_6) : $signed(_GEN_527); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_529 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_6) : $signed(_GEN_528); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_530 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_6) : $signed(_GEN_529); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_531 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_6) : $signed(_GEN_530); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_532 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_6) : $signed(_GEN_531); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_533 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_6) : $signed(_GEN_532); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_534 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_6) : $signed(_GEN_533); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_535 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_6) : $signed(_GEN_534); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_536 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_6) : $signed(_GEN_535); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_537 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_6) : $signed(_GEN_536); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_538 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_6) : $signed(_GEN_537); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_539 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_6) : $signed(_GEN_538); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_540 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_6) : $signed(_GEN_539); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_541 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_6) : $signed(_GEN_540); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_542 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_6) : $signed(_GEN_541); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_543 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_6) : $signed(_GEN_542); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_544 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_6) : $signed(_GEN_543); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_545 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_6) : $signed(_GEN_544); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_546 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_6) : $signed(_GEN_545); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_547 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_6) : $signed(_GEN_546); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_548 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_6) : $signed(_GEN_547); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_549 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_6) : $signed(_GEN_548); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_550 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_6) : $signed(_GEN_549); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_551 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_6) : $signed(_GEN_550); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_552 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_6) : $signed(_GEN_551); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_553 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_6) : $signed(_GEN_552); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_554 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_6) : $signed(_GEN_553); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_555 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_6) : $signed(_GEN_554); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_556 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_6) : $signed(_GEN_555); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_557 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_6) : $signed(_GEN_556); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_558 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_6) : $signed(_GEN_557); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_559 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_6) : $signed(_GEN_558); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_560 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_6) : $signed(_GEN_559); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_561 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_6) : $signed(_GEN_560); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_562 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_6) : $signed(_GEN_561); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_563 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_6) : $signed(_GEN_562); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_564 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_6) : $signed(_GEN_563); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_565 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_6) : $signed(_GEN_564); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_566 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_6) : $signed(_GEN_565); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_567 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_6) : $signed(_GEN_566); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_568 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_6) : $signed(_GEN_567); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_569 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_6) : $signed(_GEN_568); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_570 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_6) : $signed(_GEN_569); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_571 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_6) : $signed(_GEN_570); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_572 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_6) : $signed(_GEN_571); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_573 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_6) : $signed(_GEN_572); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_574 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_6) : $signed(_GEN_573); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_575 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_6) : $signed(_GEN_574); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_576 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_6) : $signed(_GEN_575); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_577 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_6) : $signed(_GEN_576); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_578 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_6) : $signed(_GEN_577); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_579 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_6) : $signed(_GEN_578); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_580 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_6) : $signed(_GEN_579); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_581 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_6) : $signed(_GEN_580); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_582 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_6) : $signed(_GEN_581); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_583 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_6) : $signed(_GEN_582); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_584 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_6) : $signed(_GEN_583); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_585 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_6) : $signed(_GEN_584); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_587 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_7) : $signed(cache_0_7); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_588 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_7) : $signed(_GEN_587); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_589 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_7) : $signed(_GEN_588); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_590 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_7) : $signed(_GEN_589); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_591 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_7) : $signed(_GEN_590); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_592 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_7) : $signed(_GEN_591); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_593 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_7) : $signed(_GEN_592); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_594 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_7) : $signed(_GEN_593); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_595 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_7) : $signed(_GEN_594); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_596 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_7) : $signed(_GEN_595); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_597 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_7) : $signed(_GEN_596); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_598 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_7) : $signed(_GEN_597); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_599 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_7) : $signed(_GEN_598); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_600 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_7) : $signed(_GEN_599); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_601 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_7) : $signed(_GEN_600); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_602 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_7) : $signed(_GEN_601); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_603 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_7) : $signed(_GEN_602); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_604 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_7) : $signed(_GEN_603); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_605 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_7) : $signed(_GEN_604); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_606 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_7) : $signed(_GEN_605); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_607 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_7) : $signed(_GEN_606); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_608 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_7) : $signed(_GEN_607); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_609 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_7) : $signed(_GEN_608); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_610 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_7) : $signed(_GEN_609); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_611 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_7) : $signed(_GEN_610); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_612 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_7) : $signed(_GEN_611); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_613 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_7) : $signed(_GEN_612); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_614 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_7) : $signed(_GEN_613); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_615 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_7) : $signed(_GEN_614); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_616 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_7) : $signed(_GEN_615); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_617 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_7) : $signed(_GEN_616); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_618 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_7) : $signed(_GEN_617); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_619 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_7) : $signed(_GEN_618); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_620 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_7) : $signed(_GEN_619); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_621 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_7) : $signed(_GEN_620); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_622 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_7) : $signed(_GEN_621); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_623 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_7) : $signed(_GEN_622); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_624 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_7) : $signed(_GEN_623); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_625 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_7) : $signed(_GEN_624); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_626 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_7) : $signed(_GEN_625); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_627 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_7) : $signed(_GEN_626); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_628 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_7) : $signed(_GEN_627); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_629 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_7) : $signed(_GEN_628); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_630 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_7) : $signed(_GEN_629); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_631 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_7) : $signed(_GEN_630); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_632 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_7) : $signed(_GEN_631); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_633 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_7) : $signed(_GEN_632); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_634 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_7) : $signed(_GEN_633); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_635 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_7) : $signed(_GEN_634); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_636 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_7) : $signed(_GEN_635); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_637 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_7) : $signed(_GEN_636); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_638 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_7) : $signed(_GEN_637); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_639 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_7) : $signed(_GEN_638); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_640 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_7) : $signed(_GEN_639); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_641 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_7) : $signed(_GEN_640); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_642 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_7) : $signed(_GEN_641); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_643 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_7) : $signed(_GEN_642); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_644 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_7) : $signed(_GEN_643); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_645 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_7) : $signed(_GEN_644); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_646 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_7) : $signed(_GEN_645); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_647 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_7) : $signed(_GEN_646); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_648 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_7) : $signed(_GEN_647); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_649 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_7) : $signed(_GEN_648); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_651 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_8) : $signed(cache_0_8); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_652 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_8) : $signed(_GEN_651); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_653 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_8) : $signed(_GEN_652); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_654 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_8) : $signed(_GEN_653); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_655 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_8) : $signed(_GEN_654); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_656 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_8) : $signed(_GEN_655); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_657 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_8) : $signed(_GEN_656); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_658 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_8) : $signed(_GEN_657); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_659 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_8) : $signed(_GEN_658); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_660 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_8) : $signed(_GEN_659); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_661 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_8) : $signed(_GEN_660); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_662 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_8) : $signed(_GEN_661); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_663 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_8) : $signed(_GEN_662); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_664 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_8) : $signed(_GEN_663); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_665 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_8) : $signed(_GEN_664); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_666 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_8) : $signed(_GEN_665); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_667 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_8) : $signed(_GEN_666); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_668 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_8) : $signed(_GEN_667); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_669 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_8) : $signed(_GEN_668); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_670 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_8) : $signed(_GEN_669); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_671 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_8) : $signed(_GEN_670); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_672 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_8) : $signed(_GEN_671); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_673 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_8) : $signed(_GEN_672); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_674 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_8) : $signed(_GEN_673); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_675 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_8) : $signed(_GEN_674); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_676 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_8) : $signed(_GEN_675); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_677 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_8) : $signed(_GEN_676); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_678 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_8) : $signed(_GEN_677); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_679 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_8) : $signed(_GEN_678); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_680 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_8) : $signed(_GEN_679); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_681 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_8) : $signed(_GEN_680); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_682 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_8) : $signed(_GEN_681); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_683 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_8) : $signed(_GEN_682); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_684 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_8) : $signed(_GEN_683); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_685 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_8) : $signed(_GEN_684); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_686 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_8) : $signed(_GEN_685); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_687 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_8) : $signed(_GEN_686); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_688 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_8) : $signed(_GEN_687); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_689 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_8) : $signed(_GEN_688); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_690 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_8) : $signed(_GEN_689); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_691 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_8) : $signed(_GEN_690); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_692 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_8) : $signed(_GEN_691); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_693 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_8) : $signed(_GEN_692); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_694 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_8) : $signed(_GEN_693); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_695 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_8) : $signed(_GEN_694); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_696 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_8) : $signed(_GEN_695); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_697 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_8) : $signed(_GEN_696); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_698 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_8) : $signed(_GEN_697); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_699 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_8) : $signed(_GEN_698); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_700 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_8) : $signed(_GEN_699); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_701 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_8) : $signed(_GEN_700); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_702 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_8) : $signed(_GEN_701); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_703 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_8) : $signed(_GEN_702); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_704 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_8) : $signed(_GEN_703); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_705 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_8) : $signed(_GEN_704); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_706 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_8) : $signed(_GEN_705); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_707 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_8) : $signed(_GEN_706); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_708 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_8) : $signed(_GEN_707); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_709 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_8) : $signed(_GEN_708); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_710 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_8) : $signed(_GEN_709); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_711 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_8) : $signed(_GEN_710); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_712 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_8) : $signed(_GEN_711); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_713 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_8) : $signed(_GEN_712); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_715 = 6'h1 == cnt_ic_ccnt[5:0] ? $signed(cache_1_9) : $signed(cache_0_9); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_716 = 6'h2 == cnt_ic_ccnt[5:0] ? $signed(cache_2_9) : $signed(_GEN_715); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_717 = 6'h3 == cnt_ic_ccnt[5:0] ? $signed(cache_3_9) : $signed(_GEN_716); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_718 = 6'h4 == cnt_ic_ccnt[5:0] ? $signed(cache_4_9) : $signed(_GEN_717); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_719 = 6'h5 == cnt_ic_ccnt[5:0] ? $signed(cache_5_9) : $signed(_GEN_718); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_720 = 6'h6 == cnt_ic_ccnt[5:0] ? $signed(cache_6_9) : $signed(_GEN_719); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_721 = 6'h7 == cnt_ic_ccnt[5:0] ? $signed(cache_7_9) : $signed(_GEN_720); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_722 = 6'h8 == cnt_ic_ccnt[5:0] ? $signed(cache_8_9) : $signed(_GEN_721); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_723 = 6'h9 == cnt_ic_ccnt[5:0] ? $signed(cache_9_9) : $signed(_GEN_722); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_724 = 6'ha == cnt_ic_ccnt[5:0] ? $signed(cache_10_9) : $signed(_GEN_723); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_725 = 6'hb == cnt_ic_ccnt[5:0] ? $signed(cache_11_9) : $signed(_GEN_724); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_726 = 6'hc == cnt_ic_ccnt[5:0] ? $signed(cache_12_9) : $signed(_GEN_725); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_727 = 6'hd == cnt_ic_ccnt[5:0] ? $signed(cache_13_9) : $signed(_GEN_726); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_728 = 6'he == cnt_ic_ccnt[5:0] ? $signed(cache_14_9) : $signed(_GEN_727); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_729 = 6'hf == cnt_ic_ccnt[5:0] ? $signed(cache_15_9) : $signed(_GEN_728); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_730 = 6'h10 == cnt_ic_ccnt[5:0] ? $signed(cache_16_9) : $signed(_GEN_729); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_731 = 6'h11 == cnt_ic_ccnt[5:0] ? $signed(cache_17_9) : $signed(_GEN_730); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_732 = 6'h12 == cnt_ic_ccnt[5:0] ? $signed(cache_18_9) : $signed(_GEN_731); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_733 = 6'h13 == cnt_ic_ccnt[5:0] ? $signed(cache_19_9) : $signed(_GEN_732); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_734 = 6'h14 == cnt_ic_ccnt[5:0] ? $signed(cache_20_9) : $signed(_GEN_733); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_735 = 6'h15 == cnt_ic_ccnt[5:0] ? $signed(cache_21_9) : $signed(_GEN_734); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_736 = 6'h16 == cnt_ic_ccnt[5:0] ? $signed(cache_22_9) : $signed(_GEN_735); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_737 = 6'h17 == cnt_ic_ccnt[5:0] ? $signed(cache_23_9) : $signed(_GEN_736); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_738 = 6'h18 == cnt_ic_ccnt[5:0] ? $signed(cache_24_9) : $signed(_GEN_737); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_739 = 6'h19 == cnt_ic_ccnt[5:0] ? $signed(cache_25_9) : $signed(_GEN_738); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_740 = 6'h1a == cnt_ic_ccnt[5:0] ? $signed(cache_26_9) : $signed(_GEN_739); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_741 = 6'h1b == cnt_ic_ccnt[5:0] ? $signed(cache_27_9) : $signed(_GEN_740); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_742 = 6'h1c == cnt_ic_ccnt[5:0] ? $signed(cache_28_9) : $signed(_GEN_741); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_743 = 6'h1d == cnt_ic_ccnt[5:0] ? $signed(cache_29_9) : $signed(_GEN_742); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_744 = 6'h1e == cnt_ic_ccnt[5:0] ? $signed(cache_30_9) : $signed(_GEN_743); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_745 = 6'h1f == cnt_ic_ccnt[5:0] ? $signed(cache_31_9) : $signed(_GEN_744); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_746 = 6'h20 == cnt_ic_ccnt[5:0] ? $signed(cache_32_9) : $signed(_GEN_745); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_747 = 6'h21 == cnt_ic_ccnt[5:0] ? $signed(cache_33_9) : $signed(_GEN_746); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_748 = 6'h22 == cnt_ic_ccnt[5:0] ? $signed(cache_34_9) : $signed(_GEN_747); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_749 = 6'h23 == cnt_ic_ccnt[5:0] ? $signed(cache_35_9) : $signed(_GEN_748); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_750 = 6'h24 == cnt_ic_ccnt[5:0] ? $signed(cache_36_9) : $signed(_GEN_749); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_751 = 6'h25 == cnt_ic_ccnt[5:0] ? $signed(cache_37_9) : $signed(_GEN_750); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_752 = 6'h26 == cnt_ic_ccnt[5:0] ? $signed(cache_38_9) : $signed(_GEN_751); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_753 = 6'h27 == cnt_ic_ccnt[5:0] ? $signed(cache_39_9) : $signed(_GEN_752); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_754 = 6'h28 == cnt_ic_ccnt[5:0] ? $signed(cache_40_9) : $signed(_GEN_753); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_755 = 6'h29 == cnt_ic_ccnt[5:0] ? $signed(cache_41_9) : $signed(_GEN_754); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_756 = 6'h2a == cnt_ic_ccnt[5:0] ? $signed(cache_42_9) : $signed(_GEN_755); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_757 = 6'h2b == cnt_ic_ccnt[5:0] ? $signed(cache_43_9) : $signed(_GEN_756); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_758 = 6'h2c == cnt_ic_ccnt[5:0] ? $signed(cache_44_9) : $signed(_GEN_757); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_759 = 6'h2d == cnt_ic_ccnt[5:0] ? $signed(cache_45_9) : $signed(_GEN_758); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_760 = 6'h2e == cnt_ic_ccnt[5:0] ? $signed(cache_46_9) : $signed(_GEN_759); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_761 = 6'h2f == cnt_ic_ccnt[5:0] ? $signed(cache_47_9) : $signed(_GEN_760); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_762 = 6'h30 == cnt_ic_ccnt[5:0] ? $signed(cache_48_9) : $signed(_GEN_761); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_763 = 6'h31 == cnt_ic_ccnt[5:0] ? $signed(cache_49_9) : $signed(_GEN_762); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_764 = 6'h32 == cnt_ic_ccnt[5:0] ? $signed(cache_50_9) : $signed(_GEN_763); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_765 = 6'h33 == cnt_ic_ccnt[5:0] ? $signed(cache_51_9) : $signed(_GEN_764); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_766 = 6'h34 == cnt_ic_ccnt[5:0] ? $signed(cache_52_9) : $signed(_GEN_765); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_767 = 6'h35 == cnt_ic_ccnt[5:0] ? $signed(cache_53_9) : $signed(_GEN_766); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_768 = 6'h36 == cnt_ic_ccnt[5:0] ? $signed(cache_54_9) : $signed(_GEN_767); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_769 = 6'h37 == cnt_ic_ccnt[5:0] ? $signed(cache_55_9) : $signed(_GEN_768); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_770 = 6'h38 == cnt_ic_ccnt[5:0] ? $signed(cache_56_9) : $signed(_GEN_769); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_771 = 6'h39 == cnt_ic_ccnt[5:0] ? $signed(cache_57_9) : $signed(_GEN_770); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_772 = 6'h3a == cnt_ic_ccnt[5:0] ? $signed(cache_58_9) : $signed(_GEN_771); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_773 = 6'h3b == cnt_ic_ccnt[5:0] ? $signed(cache_59_9) : $signed(_GEN_772); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_774 = 6'h3c == cnt_ic_ccnt[5:0] ? $signed(cache_60_9) : $signed(_GEN_773); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_775 = 6'h3d == cnt_ic_ccnt[5:0] ? $signed(cache_61_9) : $signed(_GEN_774); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_776 = 6'h3e == cnt_ic_ccnt[5:0] ? $signed(cache_62_9) : $signed(_GEN_775); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_777 = 6'h3f == cnt_ic_ccnt[5:0] ? $signed(cache_63_9) : $signed(_GEN_776); // @[read_pack.scala 73:26 read_pack.scala 73:26]
  wire [15:0] _GEN_778 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_21) : $signed(_GEN_329); // @[read_pack.scala 57:31 read_pack.scala 59:33 read_pack.scala 73:26]
  wire [15:0] _GEN_779 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_23) : $signed(_GEN_393); // @[read_pack.scala 57:31 read_pack.scala 59:33 read_pack.scala 73:26]
  wire [15:0] _GEN_780 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_25) : $signed(_GEN_457); // @[read_pack.scala 57:31 read_pack.scala 59:33 read_pack.scala 73:26]
  wire [15:0] _GEN_781 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_27) : $signed(_GEN_521); // @[read_pack.scala 57:31 read_pack.scala 59:33 read_pack.scala 73:26]
  wire [15:0] _GEN_782 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_29) : $signed(_GEN_585); // @[read_pack.scala 57:31 read_pack.scala 59:33 read_pack.scala 73:26]
  wire [15:0] _GEN_783 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_31) : $signed(_GEN_649); // @[read_pack.scala 57:31 read_pack.scala 59:33 read_pack.scala 73:26]
  wire [15:0] _GEN_784 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_33) : $signed(_GEN_265); // @[read_pack.scala 57:31 read_pack.scala 60:29 read_pack.scala 73:26]
  wire [15:0] _GEN_785 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_35) : $signed(_GEN_713); // @[read_pack.scala 57:31 read_pack.scala 61:29 read_pack.scala 73:26]
  wire [15:0] _GEN_786 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_134) : $signed(_GEN_201); // @[read_pack.scala 57:31 read_pack.scala 73:26]
  wire [15:0] _GEN_787 = cnt_y_ccnt == 10'h0 ? $signed(_GEN_137) : $signed(_GEN_777); // @[read_pack.scala 57:31 read_pack.scala 73:26]
  wire [15:0] _GEN_789 = state ? $signed(io_from_small_1_0_data_6) : $signed(io_from_small_0_0_data_6); // @[read_pack.scala 84:35 read_pack.scala 84:35]
  wire [15:0] _GEN_790 = _T_1 ? $signed(_GEN_101) : $signed(_GEN_789); // @[read_pack.scala 81:35 read_pack.scala 82:35 read_pack.scala 84:35]
  wire [15:0] _GEN_792 = state ? $signed(io_from_small_1_3_data_6) : $signed(io_from_small_0_3_data_6); // @[read_pack.scala 89:35 read_pack.scala 89:35]
  wire [15:0] _GEN_793 = nxt_2 ? $signed(_GEN_111) : $signed(_GEN_792); // @[read_pack.scala 86:42 read_pack.scala 87:35 read_pack.scala 89:35]
  wire [15:0] _GEN_795 = _state_T ? $signed(io_from_big_1_data_0) : $signed(io_from_big_0_data_0); // @[read_pack.scala 93:35 read_pack.scala 93:35]
  wire [15:0] _GEN_797 = _state_T ? $signed(io_from_big_1_data_1) : $signed(io_from_big_0_data_1); // @[read_pack.scala 93:35 read_pack.scala 93:35]
  wire [15:0] _GEN_799 = _state_T ? $signed(io_from_big_1_data_2) : $signed(io_from_big_0_data_2); // @[read_pack.scala 93:35 read_pack.scala 93:35]
  wire [15:0] _GEN_801 = _state_T ? $signed(io_from_big_1_data_3) : $signed(io_from_big_0_data_3); // @[read_pack.scala 93:35 read_pack.scala 93:35]
  wire [15:0] _GEN_803 = _state_T ? $signed(io_from_big_1_data_4) : $signed(io_from_big_0_data_4); // @[read_pack.scala 93:35 read_pack.scala 93:35]
  wire [15:0] _GEN_805 = _state_T ? $signed(io_from_big_1_data_5) : $signed(io_from_big_0_data_5); // @[read_pack.scala 93:35 read_pack.scala 93:35]
  wire [15:0] _GEN_807 = _state_T ? $signed(io_from_small_1_1_data_0) : $signed(io_from_small_0_1_data_0); // @[read_pack.scala 94:31 read_pack.scala 94:31]
  wire [15:0] _GEN_809 = _state_T ? $signed(io_from_small_1_2_data_0) : $signed(io_from_small_0_2_data_0); // @[read_pack.scala 95:31 read_pack.scala 95:31]
  wire [15:0] _GEN_813 = _state_T ? $signed(io_from_small_1_0_data_0) : $signed(io_from_small_0_0_data_0); // @[read_pack.scala 99:35 read_pack.scala 99:35]
  wire [15:0] _GEN_814 = _T_1 ? $signed(_GEN_795) : $signed(_GEN_813); // @[read_pack.scala 96:35 read_pack.scala 97:35 read_pack.scala 99:35]
  wire [15:0] _GEN_818 = _state_T ? $signed(io_from_small_1_3_data_0) : $signed(io_from_small_0_3_data_0); // @[read_pack.scala 104:35 read_pack.scala 104:35]
  wire [15:0] _GEN_819 = nxt_2 ? $signed(_GEN_805) : $signed(_GEN_818); // @[read_pack.scala 101:42 read_pack.scala 102:35 read_pack.scala 104:35]
  wire [15:0] _GEN_820 = nxt_1 ? $signed(_GEN_101) : $signed(_GEN_795); // @[read_pack.scala 76:38 read_pack.scala 78:35 read_pack.scala 93:35]
  wire [15:0] _GEN_821 = nxt_1 ? $signed(_GEN_103) : $signed(_GEN_797); // @[read_pack.scala 76:38 read_pack.scala 78:35 read_pack.scala 93:35]
  wire [15:0] _GEN_822 = nxt_1 ? $signed(_GEN_105) : $signed(_GEN_799); // @[read_pack.scala 76:38 read_pack.scala 78:35 read_pack.scala 93:35]
  wire [15:0] _GEN_823 = nxt_1 ? $signed(_GEN_107) : $signed(_GEN_801); // @[read_pack.scala 76:38 read_pack.scala 78:35 read_pack.scala 93:35]
  wire [15:0] _GEN_824 = nxt_1 ? $signed(_GEN_109) : $signed(_GEN_803); // @[read_pack.scala 76:38 read_pack.scala 78:35 read_pack.scala 93:35]
  wire [15:0] _GEN_825 = nxt_1 ? $signed(_GEN_111) : $signed(_GEN_805); // @[read_pack.scala 76:38 read_pack.scala 78:35 read_pack.scala 93:35]
  wire [15:0] _GEN_826 = nxt_1 ? $signed(_GEN_113) : $signed(_GEN_807); // @[read_pack.scala 76:38 read_pack.scala 79:31 read_pack.scala 94:31]
  wire [15:0] _GEN_827 = nxt_1 ? $signed(_GEN_115) : $signed(_GEN_809); // @[read_pack.scala 76:38 read_pack.scala 80:31 read_pack.scala 95:31]
  wire [15:0] _GEN_828 = nxt_1 ? $signed(_GEN_790) : $signed(_GEN_814); // @[read_pack.scala 76:38]
  wire [15:0] _GEN_829 = nxt_1 ? $signed(_GEN_793) : $signed(_GEN_819); // @[read_pack.scala 76:38]
  wire [15:0] _GEN_831 = state ? $signed(io_from_small_1_0_data_0) : $signed(io_from_small_0_0_data_0); // @[read_pack.scala 112:28 read_pack.scala 112:28]
  wire [15:0] _GEN_833 = state ? $signed(io_from_small_1_0_data_2) : $signed(io_from_small_0_0_data_2); // @[read_pack.scala 112:28 read_pack.scala 112:28]
  wire [15:0] _GEN_835 = state ? $signed(io_from_small_1_0_data_3) : $signed(io_from_small_0_0_data_3); // @[read_pack.scala 112:28 read_pack.scala 112:28]
  wire [15:0] _GEN_837 = state ? $signed(io_from_small_1_0_data_4) : $signed(io_from_small_0_0_data_4); // @[read_pack.scala 112:28 read_pack.scala 112:28]
  wire [15:0] _GEN_839 = state ? $signed(io_from_small_1_0_data_5) : $signed(io_from_small_0_0_data_5); // @[read_pack.scala 112:28 read_pack.scala 112:28]
  wire [15:0] _GEN_841 = state ? $signed(io_from_small_1_0_data_7) : $signed(io_from_small_0_0_data_7); // @[read_pack.scala 112:28 read_pack.scala 112:28]
  wire [15:0] _GEN_842 = _T_1 ? $signed(_GEN_5) : $signed(_GEN_831); // @[read_pack.scala 108:31 read_pack.scala 110:35 read_pack.scala 112:28]
  wire [15:0] _GEN_844 = _T_1 ? $signed(_GEN_37) : $signed(_GEN_833); // @[read_pack.scala 108:31 read_pack.scala 110:35 read_pack.scala 112:28]
  wire [15:0] _GEN_845 = _T_1 ? $signed(_GEN_53) : $signed(_GEN_835); // @[read_pack.scala 108:31 read_pack.scala 110:35 read_pack.scala 112:28]
  wire [15:0] _GEN_846 = _T_1 ? $signed(_GEN_69) : $signed(_GEN_837); // @[read_pack.scala 108:31 read_pack.scala 110:35 read_pack.scala 112:28]
  wire [15:0] _GEN_847 = _T_1 ? $signed(_GEN_85) : $signed(_GEN_839); // @[read_pack.scala 108:31 read_pack.scala 110:35 read_pack.scala 112:28]
  wire [15:0] _GEN_849 = _T_1 ? $signed(nxt_up_2) : $signed(_GEN_841); // @[read_pack.scala 108:31 read_pack.scala 110:35 read_pack.scala 112:28]
  wire [15:0] _GEN_851 = state ? $signed(io_from_small_1_3_data_0) : $signed(io_from_small_0_3_data_0); // @[read_pack.scala 118:29 read_pack.scala 118:29]
  wire [15:0] _GEN_853 = state ? $signed(io_from_small_1_3_data_2) : $signed(io_from_small_0_3_data_2); // @[read_pack.scala 118:29 read_pack.scala 118:29]
  wire [15:0] _GEN_855 = state ? $signed(io_from_small_1_3_data_3) : $signed(io_from_small_0_3_data_3); // @[read_pack.scala 118:29 read_pack.scala 118:29]
  wire [15:0] _GEN_857 = state ? $signed(io_from_small_1_3_data_4) : $signed(io_from_small_0_3_data_4); // @[read_pack.scala 118:29 read_pack.scala 118:29]
  wire [15:0] _GEN_859 = state ? $signed(io_from_small_1_3_data_5) : $signed(io_from_small_0_3_data_5); // @[read_pack.scala 118:29 read_pack.scala 118:29]
  wire [15:0] _GEN_861 = state ? $signed(io_from_small_1_3_data_7) : $signed(io_from_small_0_3_data_7); // @[read_pack.scala 118:29 read_pack.scala 118:29]
  wire [15:0] _GEN_862 = nxt_2 ? $signed(_GEN_15) : $signed(_GEN_851); // @[read_pack.scala 114:38 read_pack.scala 116:36 read_pack.scala 118:29]
  wire [15:0] _GEN_864 = nxt_2 ? $signed(_GEN_47) : $signed(_GEN_853); // @[read_pack.scala 114:38 read_pack.scala 116:36 read_pack.scala 118:29]
  wire [15:0] _GEN_865 = nxt_2 ? $signed(_GEN_63) : $signed(_GEN_855); // @[read_pack.scala 114:38 read_pack.scala 116:36 read_pack.scala 118:29]
  wire [15:0] _GEN_866 = nxt_2 ? $signed(_GEN_79) : $signed(_GEN_857); // @[read_pack.scala 114:38 read_pack.scala 116:36 read_pack.scala 118:29]
  wire [15:0] _GEN_867 = nxt_2 ? $signed(_GEN_95) : $signed(_GEN_859); // @[read_pack.scala 114:38 read_pack.scala 116:36 read_pack.scala 118:29]
  wire [15:0] _GEN_869 = nxt_2 ? $signed(nxt_up_7) : $signed(_GEN_861); // @[read_pack.scala 114:38 read_pack.scala 116:36 read_pack.scala 118:29]
  wire [15:0] _GEN_1517 = io_valid_in ? $signed(_GEN_5) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1518 = io_valid_in ? $signed(_GEN_7) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1519 = io_valid_in ? $signed(_GEN_9) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1520 = io_valid_in ? $signed(_GEN_11) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1521 = io_valid_in ? $signed(_GEN_13) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1522 = io_valid_in ? $signed(_GEN_15) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1523 = io_valid_in ? $signed(_GEN_17) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 39:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1524 = io_valid_in ? $signed(_GEN_19) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 40:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1525 = io_valid_in ? $signed(_GEN_21) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1526 = io_valid_in ? $signed(_GEN_23) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1527 = io_valid_in ? $signed(_GEN_25) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1528 = io_valid_in ? $signed(_GEN_27) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1529 = io_valid_in ? $signed(_GEN_29) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1530 = io_valid_in ? $signed(_GEN_31) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1531 = io_valid_in ? $signed(_GEN_33) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 39:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1532 = io_valid_in ? $signed(_GEN_35) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 40:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1533 = io_valid_in ? $signed(_GEN_37) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1534 = io_valid_in ? $signed(_GEN_39) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1535 = io_valid_in ? $signed(_GEN_41) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1536 = io_valid_in ? $signed(_GEN_43) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1537 = io_valid_in ? $signed(_GEN_45) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1538 = io_valid_in ? $signed(_GEN_47) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1539 = io_valid_in ? $signed(_GEN_49) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 39:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1540 = io_valid_in ? $signed(_GEN_51) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 40:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1541 = io_valid_in ? $signed(_GEN_53) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1542 = io_valid_in ? $signed(_GEN_55) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1543 = io_valid_in ? $signed(_GEN_57) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1544 = io_valid_in ? $signed(_GEN_59) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1545 = io_valid_in ? $signed(_GEN_61) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1546 = io_valid_in ? $signed(_GEN_63) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1547 = io_valid_in ? $signed(_GEN_65) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 39:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1548 = io_valid_in ? $signed(_GEN_67) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 40:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1549 = io_valid_in ? $signed(_GEN_69) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1550 = io_valid_in ? $signed(_GEN_71) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1551 = io_valid_in ? $signed(_GEN_73) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1552 = io_valid_in ? $signed(_GEN_75) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1553 = io_valid_in ? $signed(_GEN_77) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1554 = io_valid_in ? $signed(_GEN_79) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1555 = io_valid_in ? $signed(_GEN_81) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 39:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1556 = io_valid_in ? $signed(_GEN_83) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 40:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1557 = io_valid_in ? $signed(_GEN_85) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1558 = io_valid_in ? $signed(_GEN_87) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1559 = io_valid_in ? $signed(_GEN_89) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1560 = io_valid_in ? $signed(_GEN_91) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1561 = io_valid_in ? $signed(_GEN_93) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1562 = io_valid_in ? $signed(_GEN_95) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1563 = io_valid_in ? $signed(_GEN_97) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 39:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1564 = io_valid_in ? $signed(_GEN_99) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 40:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1565 = io_valid_in ? $signed(_GEN_101) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1566 = io_valid_in ? $signed(_GEN_103) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1567 = io_valid_in ? $signed(_GEN_105) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1568 = io_valid_in ? $signed(_GEN_107) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1569 = io_valid_in ? $signed(_GEN_109) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1570 = io_valid_in ? $signed(_GEN_111) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1571 = io_valid_in ? $signed(_GEN_113) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 39:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1572 = io_valid_in ? $signed(_GEN_115) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 40:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1573 = io_valid_in ? $signed(nxt_up_2) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1574 = io_valid_in ? $signed(nxt_up_3) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1575 = io_valid_in ? $signed(nxt_up_4) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1576 = io_valid_in ? $signed(nxt_up_5) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1577 = io_valid_in ? $signed(nxt_up_6) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1578 = io_valid_in ? $signed(nxt_up_7) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 38:38 read_pack.scala 30:15]
  wire [15:0] _GEN_1579 = io_valid_in ? $signed(nxt_up_1) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 39:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1580 = io_valid_in ? $signed(nxt_up_8) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 40:34 read_pack.scala 30:15]
  wire [15:0] _GEN_1581 = io_valid_in ? $signed(_GEN_778) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1582 = io_valid_in ? $signed(_GEN_779) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1583 = io_valid_in ? $signed(_GEN_780) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1584 = io_valid_in ? $signed(_GEN_781) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1585 = io_valid_in ? $signed(_GEN_782) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1586 = io_valid_in ? $signed(_GEN_783) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1587 = io_valid_in ? $signed(_GEN_784) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1588 = io_valid_in ? $signed(_GEN_785) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1589 = io_valid_in ? $signed(_GEN_786) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1590 = io_valid_in ? $signed(_GEN_787) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1591 = io_valid_in ? $signed(_GEN_820) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1592 = io_valid_in ? $signed(_GEN_821) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1593 = io_valid_in ? $signed(_GEN_822) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1594 = io_valid_in ? $signed(_GEN_823) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1595 = io_valid_in ? $signed(_GEN_824) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1596 = io_valid_in ? $signed(_GEN_825) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1597 = io_valid_in ? $signed(_GEN_826) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1598 = io_valid_in ? $signed(_GEN_827) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1599 = io_valid_in ? $signed(_GEN_828) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1600 = io_valid_in ? $signed(_GEN_829) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1601 = io_valid_in ? $signed(_GEN_842) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1602 = io_valid_in ? $signed(_GEN_134) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1603 = io_valid_in ? $signed(_GEN_844) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1604 = io_valid_in ? $signed(_GEN_845) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1605 = io_valid_in ? $signed(_GEN_846) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1606 = io_valid_in ? $signed(_GEN_847) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1607 = io_valid_in ? $signed(_GEN_790) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1608 = io_valid_in ? $signed(_GEN_849) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1609 = io_valid_in ? $signed(_GEN_862) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1610 = io_valid_in ? $signed(_GEN_137) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1611 = io_valid_in ? $signed(_GEN_864) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1612 = io_valid_in ? $signed(_GEN_865) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1613 = io_valid_in ? $signed(_GEN_866) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1614 = io_valid_in ? $signed(_GEN_867) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1615 = io_valid_in ? $signed(_GEN_793) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  wire [15:0] _GEN_1616 = io_valid_in ? $signed(_GEN_869) : $signed(16'sh0); // @[read_pack.scala 48:28 read_pack.scala 30:15]
  assign io_valid_out = io_flag_job ? 1'h0 : io_valid_in; // @[read_pack.scala 43:22 read_pack.scala 29:18]
  assign io_output_mat_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1523); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1517); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1518); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1519); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1520); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1521); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1522); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1524); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1531); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1525); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_10 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1526); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_11 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1527); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_12 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1528); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_13 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1529); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_14 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1530); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_15 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1532); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_16 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1539); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_17 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1533); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_18 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1534); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_19 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1535); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_20 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1536); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_21 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1537); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_22 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1538); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_23 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1540); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_24 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1547); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_25 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1541); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_26 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1542); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_27 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1543); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_28 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1544); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_29 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1545); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_30 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1546); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_31 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1548); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_32 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1555); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_33 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1549); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_34 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1550); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_35 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1551); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_36 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1552); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_37 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1553); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_38 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1554); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_39 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1556); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_40 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1563); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_41 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1557); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_42 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1558); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_43 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1559); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_44 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1560); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_45 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1561); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_46 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1562); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_47 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1564); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_48 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1571); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_49 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1565); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_50 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1566); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_51 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1567); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_52 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1568); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_53 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1569); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_54 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1570); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_55 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1572); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_56 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1579); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_57 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1573); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_58 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1574); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_59 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1575); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_60 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1576); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_61 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1577); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_62 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1578); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_mat_63 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1580); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1589); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1587); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1581); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1582); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1583); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1584); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1585); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1586); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1588); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_up_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1590); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1599); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1597); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1591); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1592); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1593); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1594); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1595); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1596); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1598); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_down_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1600); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_left_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1601); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_left_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1602); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_left_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1603); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_left_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1604); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_left_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1605); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_left_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1606); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_left_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1607); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_left_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1608); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_right_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1609); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_right_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1610); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_right_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1611); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_right_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1612); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_right_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1613); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_right_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1614); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_right_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1615); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  assign io_output_right_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1616); // @[read_pack.scala 43:22 read_pack.scala 30:15]
  always @(posedge clock) begin
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_0_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h0 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_0_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_1_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_1_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_2_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_2_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_3_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_3_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_4_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h4 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_4_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_5_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h5 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_5_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_6_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h6 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_6_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_7_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h7 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_7_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_8_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h8 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_8_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_9_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h9 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_9_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_10_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'ha == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_10_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_11_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hb == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_11_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_12_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hc == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_12_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_13_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hd == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_13_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_14_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'he == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_14_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_15_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'hf == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_15_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_16_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h10 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_16_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_17_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h11 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_17_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_18_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h12 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_18_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_19_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h13 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_19_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_20_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h14 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_20_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_21_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h15 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_21_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_22_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h16 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_22_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_23_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h17 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_23_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_24_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h18 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_24_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_25_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h19 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_25_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_26_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_26_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_27_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_27_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_28_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_28_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_29_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_29_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_30_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_30_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_31_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h1f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_31_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_32_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h20 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_32_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_33_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h21 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_33_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_34_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h22 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_34_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_35_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h23 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_35_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_36_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h24 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_36_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_37_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h25 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_37_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_38_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h26 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_38_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_39_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h27 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_39_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_40_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h28 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_40_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_41_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h29 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_41_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_42_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_42_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_43_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_43_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_44_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_44_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_45_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_45_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_46_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_46_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_47_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h2f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_47_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_48_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h30 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_48_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_49_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h31 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_49_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_50_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h32 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_50_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_51_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h33 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_51_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_52_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h34 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_52_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_53_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h35 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_53_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_54_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h36 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_54_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_55_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h37 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_55_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_56_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h38 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_56_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_57_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h39 == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_57_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_58_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3a == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_58_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_59_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3b == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_59_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_60_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3c == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_60_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_61_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3d == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_61_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_62_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3e == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_62_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_0 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_0 <= _GEN_849; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_1 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_1 <= nxt_up_1; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_2 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_2 <= nxt_up_2; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_3 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_3 <= nxt_up_3; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_4 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_4 <= nxt_up_4; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_5 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_5 <= nxt_up_5; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_6 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_6 <= nxt_up_6; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_7 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_7 <= nxt_up_7; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_8 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_8 <= nxt_up_8; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 23:24]
      cache_63_9 <= 16'sh0; // @[read_pack.scala 23:24]
    end else if (!(io_flag_job)) begin // @[read_pack.scala 43:22]
      if (io_valid_in) begin // @[read_pack.scala 48:28]
        if (6'h3f == cnt_ic_ccnt[5:0]) begin // @[read_pack.scala 136:28]
          cache_63_9 <= _GEN_869; // @[read_pack.scala 136:28]
        end
      end
    end
    if (reset) begin // @[read_pack.scala 25:25]
      cnt_ic_ccnt <= 10'h0; // @[read_pack.scala 25:25]
    end else if (io_flag_job) begin // @[read_pack.scala 43:22]
      cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read_pack.scala 48:28]
      if (nxt) begin // @[utils.scala 18:20]
        cnt_ic_ccnt <= 10'h0;
      end else begin
        cnt_ic_ccnt <= _cnt_ic_ccnt_T_1;
      end
    end
    if (reset) begin // @[read_pack.scala 25:25]
      cnt_ic_cend <= 10'h0; // @[read_pack.scala 25:25]
    end else if (io_flag_job) begin // @[read_pack.scala 43:22]
      cnt_ic_cend <= io_job_in_chan; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read_pack.scala 26:24]
      cnt_x_ccnt <= 10'h0; // @[read_pack.scala 26:24]
    end else if (io_flag_job) begin // @[read_pack.scala 43:22]
      cnt_x_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read_pack.scala 48:28]
      if (nxt) begin // @[read_pack.scala 50:27]
        cnt_x_ccnt <= _GEN_0;
      end
    end
    if (reset) begin // @[read_pack.scala 26:24]
      cnt_x_cend <= 10'h0; // @[read_pack.scala 26:24]
    end else if (io_flag_job) begin // @[read_pack.scala 43:22]
      cnt_x_cend <= io_job_cnt_x_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read_pack.scala 27:24]
      cnt_y_ccnt <= 10'h0; // @[read_pack.scala 27:24]
    end else if (io_flag_job) begin // @[read_pack.scala 43:22]
      cnt_y_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[read_pack.scala 48:28]
      if (nxt) begin // @[read_pack.scala 50:27]
        cnt_y_ccnt <= _cnt_y_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[read_pack.scala 27:24]
      cnt_y_cend <= 10'h0; // @[read_pack.scala 27:24]
    end else if (io_flag_job) begin // @[read_pack.scala 43:22]
      cnt_y_cend <= io_job_cnt_y_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[read_pack.scala 33:24]
      state <= 1'h0; // @[read_pack.scala 33:24]
    end else if (io_flag_job) begin // @[read_pack.scala 43:22]
      state <= 1'h0; // @[read_pack.scala 47:15]
    end else if (io_valid_in) begin // @[read_pack.scala 48:28]
      if (nxt) begin // @[read_pack.scala 50:27]
        state <= ~state; // @[read_pack.scala 51:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cache_0_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  cache_0_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  cache_0_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  cache_0_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  cache_0_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  cache_0_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  cache_0_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  cache_0_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  cache_0_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  cache_0_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  cache_1_0 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  cache_1_1 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  cache_1_2 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  cache_1_3 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  cache_1_4 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  cache_1_5 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  cache_1_6 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  cache_1_7 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  cache_1_8 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  cache_1_9 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  cache_2_0 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  cache_2_1 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  cache_2_2 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  cache_2_3 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  cache_2_4 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  cache_2_5 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  cache_2_6 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  cache_2_7 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  cache_2_8 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  cache_2_9 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  cache_3_0 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  cache_3_1 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  cache_3_2 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  cache_3_3 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  cache_3_4 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  cache_3_5 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  cache_3_6 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  cache_3_7 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  cache_3_8 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  cache_3_9 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  cache_4_0 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  cache_4_1 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  cache_4_2 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  cache_4_3 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  cache_4_4 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  cache_4_5 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  cache_4_6 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  cache_4_7 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  cache_4_8 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  cache_4_9 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  cache_5_0 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  cache_5_1 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  cache_5_2 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  cache_5_3 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  cache_5_4 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  cache_5_5 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  cache_5_6 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  cache_5_7 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  cache_5_8 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  cache_5_9 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  cache_6_0 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  cache_6_1 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  cache_6_2 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  cache_6_3 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  cache_6_4 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  cache_6_5 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  cache_6_6 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  cache_6_7 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  cache_6_8 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  cache_6_9 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  cache_7_0 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  cache_7_1 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  cache_7_2 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  cache_7_3 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  cache_7_4 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  cache_7_5 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  cache_7_6 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  cache_7_7 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  cache_7_8 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  cache_7_9 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  cache_8_0 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  cache_8_1 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  cache_8_2 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  cache_8_3 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  cache_8_4 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  cache_8_5 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  cache_8_6 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  cache_8_7 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  cache_8_8 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  cache_8_9 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  cache_9_0 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  cache_9_1 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  cache_9_2 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  cache_9_3 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  cache_9_4 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  cache_9_5 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  cache_9_6 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  cache_9_7 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  cache_9_8 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  cache_9_9 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  cache_10_0 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  cache_10_1 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  cache_10_2 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  cache_10_3 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  cache_10_4 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  cache_10_5 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  cache_10_6 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  cache_10_7 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  cache_10_8 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  cache_10_9 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  cache_11_0 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  cache_11_1 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  cache_11_2 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  cache_11_3 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  cache_11_4 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  cache_11_5 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  cache_11_6 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  cache_11_7 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  cache_11_8 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  cache_11_9 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  cache_12_0 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  cache_12_1 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  cache_12_2 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  cache_12_3 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  cache_12_4 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  cache_12_5 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  cache_12_6 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  cache_12_7 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  cache_12_8 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  cache_12_9 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  cache_13_0 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  cache_13_1 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  cache_13_2 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  cache_13_3 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  cache_13_4 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  cache_13_5 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  cache_13_6 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  cache_13_7 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  cache_13_8 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  cache_13_9 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  cache_14_0 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  cache_14_1 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  cache_14_2 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  cache_14_3 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  cache_14_4 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  cache_14_5 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  cache_14_6 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  cache_14_7 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  cache_14_8 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  cache_14_9 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  cache_15_0 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  cache_15_1 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  cache_15_2 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  cache_15_3 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  cache_15_4 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  cache_15_5 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  cache_15_6 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  cache_15_7 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  cache_15_8 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  cache_15_9 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  cache_16_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  cache_16_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  cache_16_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  cache_16_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  cache_16_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  cache_16_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  cache_16_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  cache_16_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  cache_16_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  cache_16_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  cache_17_0 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  cache_17_1 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  cache_17_2 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  cache_17_3 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  cache_17_4 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  cache_17_5 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  cache_17_6 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  cache_17_7 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  cache_17_8 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  cache_17_9 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  cache_18_0 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  cache_18_1 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  cache_18_2 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  cache_18_3 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  cache_18_4 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  cache_18_5 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  cache_18_6 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  cache_18_7 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  cache_18_8 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  cache_18_9 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  cache_19_0 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  cache_19_1 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  cache_19_2 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  cache_19_3 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  cache_19_4 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  cache_19_5 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  cache_19_6 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  cache_19_7 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  cache_19_8 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  cache_19_9 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  cache_20_0 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  cache_20_1 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  cache_20_2 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  cache_20_3 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  cache_20_4 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  cache_20_5 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  cache_20_6 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  cache_20_7 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  cache_20_8 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  cache_20_9 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  cache_21_0 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  cache_21_1 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  cache_21_2 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  cache_21_3 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  cache_21_4 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  cache_21_5 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  cache_21_6 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  cache_21_7 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  cache_21_8 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  cache_21_9 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  cache_22_0 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  cache_22_1 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  cache_22_2 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  cache_22_3 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  cache_22_4 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  cache_22_5 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  cache_22_6 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  cache_22_7 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  cache_22_8 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  cache_22_9 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  cache_23_0 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  cache_23_1 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  cache_23_2 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  cache_23_3 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  cache_23_4 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  cache_23_5 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  cache_23_6 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  cache_23_7 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  cache_23_8 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  cache_23_9 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  cache_24_0 = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  cache_24_1 = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  cache_24_2 = _RAND_242[15:0];
  _RAND_243 = {1{`RANDOM}};
  cache_24_3 = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  cache_24_4 = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  cache_24_5 = _RAND_245[15:0];
  _RAND_246 = {1{`RANDOM}};
  cache_24_6 = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  cache_24_7 = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  cache_24_8 = _RAND_248[15:0];
  _RAND_249 = {1{`RANDOM}};
  cache_24_9 = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  cache_25_0 = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  cache_25_1 = _RAND_251[15:0];
  _RAND_252 = {1{`RANDOM}};
  cache_25_2 = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  cache_25_3 = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  cache_25_4 = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  cache_25_5 = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  cache_25_6 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  cache_25_7 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  cache_25_8 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  cache_25_9 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  cache_26_0 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  cache_26_1 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  cache_26_2 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  cache_26_3 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  cache_26_4 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  cache_26_5 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  cache_26_6 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  cache_26_7 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  cache_26_8 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  cache_26_9 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  cache_27_0 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  cache_27_1 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  cache_27_2 = _RAND_272[15:0];
  _RAND_273 = {1{`RANDOM}};
  cache_27_3 = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  cache_27_4 = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  cache_27_5 = _RAND_275[15:0];
  _RAND_276 = {1{`RANDOM}};
  cache_27_6 = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  cache_27_7 = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  cache_27_8 = _RAND_278[15:0];
  _RAND_279 = {1{`RANDOM}};
  cache_27_9 = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  cache_28_0 = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  cache_28_1 = _RAND_281[15:0];
  _RAND_282 = {1{`RANDOM}};
  cache_28_2 = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  cache_28_3 = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  cache_28_4 = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  cache_28_5 = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  cache_28_6 = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  cache_28_7 = _RAND_287[15:0];
  _RAND_288 = {1{`RANDOM}};
  cache_28_8 = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  cache_28_9 = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  cache_29_0 = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  cache_29_1 = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  cache_29_2 = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  cache_29_3 = _RAND_293[15:0];
  _RAND_294 = {1{`RANDOM}};
  cache_29_4 = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  cache_29_5 = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  cache_29_6 = _RAND_296[15:0];
  _RAND_297 = {1{`RANDOM}};
  cache_29_7 = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  cache_29_8 = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  cache_29_9 = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  cache_30_0 = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  cache_30_1 = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  cache_30_2 = _RAND_302[15:0];
  _RAND_303 = {1{`RANDOM}};
  cache_30_3 = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  cache_30_4 = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  cache_30_5 = _RAND_305[15:0];
  _RAND_306 = {1{`RANDOM}};
  cache_30_6 = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  cache_30_7 = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  cache_30_8 = _RAND_308[15:0];
  _RAND_309 = {1{`RANDOM}};
  cache_30_9 = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  cache_31_0 = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  cache_31_1 = _RAND_311[15:0];
  _RAND_312 = {1{`RANDOM}};
  cache_31_2 = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  cache_31_3 = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  cache_31_4 = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  cache_31_5 = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  cache_31_6 = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  cache_31_7 = _RAND_317[15:0];
  _RAND_318 = {1{`RANDOM}};
  cache_31_8 = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  cache_31_9 = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  cache_32_0 = _RAND_320[15:0];
  _RAND_321 = {1{`RANDOM}};
  cache_32_1 = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  cache_32_2 = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  cache_32_3 = _RAND_323[15:0];
  _RAND_324 = {1{`RANDOM}};
  cache_32_4 = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  cache_32_5 = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  cache_32_6 = _RAND_326[15:0];
  _RAND_327 = {1{`RANDOM}};
  cache_32_7 = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  cache_32_8 = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  cache_32_9 = _RAND_329[15:0];
  _RAND_330 = {1{`RANDOM}};
  cache_33_0 = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  cache_33_1 = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  cache_33_2 = _RAND_332[15:0];
  _RAND_333 = {1{`RANDOM}};
  cache_33_3 = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  cache_33_4 = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  cache_33_5 = _RAND_335[15:0];
  _RAND_336 = {1{`RANDOM}};
  cache_33_6 = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  cache_33_7 = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  cache_33_8 = _RAND_338[15:0];
  _RAND_339 = {1{`RANDOM}};
  cache_33_9 = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  cache_34_0 = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  cache_34_1 = _RAND_341[15:0];
  _RAND_342 = {1{`RANDOM}};
  cache_34_2 = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  cache_34_3 = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  cache_34_4 = _RAND_344[15:0];
  _RAND_345 = {1{`RANDOM}};
  cache_34_5 = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  cache_34_6 = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  cache_34_7 = _RAND_347[15:0];
  _RAND_348 = {1{`RANDOM}};
  cache_34_8 = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  cache_34_9 = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  cache_35_0 = _RAND_350[15:0];
  _RAND_351 = {1{`RANDOM}};
  cache_35_1 = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  cache_35_2 = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  cache_35_3 = _RAND_353[15:0];
  _RAND_354 = {1{`RANDOM}};
  cache_35_4 = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  cache_35_5 = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  cache_35_6 = _RAND_356[15:0];
  _RAND_357 = {1{`RANDOM}};
  cache_35_7 = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  cache_35_8 = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  cache_35_9 = _RAND_359[15:0];
  _RAND_360 = {1{`RANDOM}};
  cache_36_0 = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  cache_36_1 = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  cache_36_2 = _RAND_362[15:0];
  _RAND_363 = {1{`RANDOM}};
  cache_36_3 = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  cache_36_4 = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  cache_36_5 = _RAND_365[15:0];
  _RAND_366 = {1{`RANDOM}};
  cache_36_6 = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  cache_36_7 = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  cache_36_8 = _RAND_368[15:0];
  _RAND_369 = {1{`RANDOM}};
  cache_36_9 = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  cache_37_0 = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  cache_37_1 = _RAND_371[15:0];
  _RAND_372 = {1{`RANDOM}};
  cache_37_2 = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  cache_37_3 = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  cache_37_4 = _RAND_374[15:0];
  _RAND_375 = {1{`RANDOM}};
  cache_37_5 = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  cache_37_6 = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  cache_37_7 = _RAND_377[15:0];
  _RAND_378 = {1{`RANDOM}};
  cache_37_8 = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  cache_37_9 = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  cache_38_0 = _RAND_380[15:0];
  _RAND_381 = {1{`RANDOM}};
  cache_38_1 = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  cache_38_2 = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  cache_38_3 = _RAND_383[15:0];
  _RAND_384 = {1{`RANDOM}};
  cache_38_4 = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  cache_38_5 = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  cache_38_6 = _RAND_386[15:0];
  _RAND_387 = {1{`RANDOM}};
  cache_38_7 = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  cache_38_8 = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  cache_38_9 = _RAND_389[15:0];
  _RAND_390 = {1{`RANDOM}};
  cache_39_0 = _RAND_390[15:0];
  _RAND_391 = {1{`RANDOM}};
  cache_39_1 = _RAND_391[15:0];
  _RAND_392 = {1{`RANDOM}};
  cache_39_2 = _RAND_392[15:0];
  _RAND_393 = {1{`RANDOM}};
  cache_39_3 = _RAND_393[15:0];
  _RAND_394 = {1{`RANDOM}};
  cache_39_4 = _RAND_394[15:0];
  _RAND_395 = {1{`RANDOM}};
  cache_39_5 = _RAND_395[15:0];
  _RAND_396 = {1{`RANDOM}};
  cache_39_6 = _RAND_396[15:0];
  _RAND_397 = {1{`RANDOM}};
  cache_39_7 = _RAND_397[15:0];
  _RAND_398 = {1{`RANDOM}};
  cache_39_8 = _RAND_398[15:0];
  _RAND_399 = {1{`RANDOM}};
  cache_39_9 = _RAND_399[15:0];
  _RAND_400 = {1{`RANDOM}};
  cache_40_0 = _RAND_400[15:0];
  _RAND_401 = {1{`RANDOM}};
  cache_40_1 = _RAND_401[15:0];
  _RAND_402 = {1{`RANDOM}};
  cache_40_2 = _RAND_402[15:0];
  _RAND_403 = {1{`RANDOM}};
  cache_40_3 = _RAND_403[15:0];
  _RAND_404 = {1{`RANDOM}};
  cache_40_4 = _RAND_404[15:0];
  _RAND_405 = {1{`RANDOM}};
  cache_40_5 = _RAND_405[15:0];
  _RAND_406 = {1{`RANDOM}};
  cache_40_6 = _RAND_406[15:0];
  _RAND_407 = {1{`RANDOM}};
  cache_40_7 = _RAND_407[15:0];
  _RAND_408 = {1{`RANDOM}};
  cache_40_8 = _RAND_408[15:0];
  _RAND_409 = {1{`RANDOM}};
  cache_40_9 = _RAND_409[15:0];
  _RAND_410 = {1{`RANDOM}};
  cache_41_0 = _RAND_410[15:0];
  _RAND_411 = {1{`RANDOM}};
  cache_41_1 = _RAND_411[15:0];
  _RAND_412 = {1{`RANDOM}};
  cache_41_2 = _RAND_412[15:0];
  _RAND_413 = {1{`RANDOM}};
  cache_41_3 = _RAND_413[15:0];
  _RAND_414 = {1{`RANDOM}};
  cache_41_4 = _RAND_414[15:0];
  _RAND_415 = {1{`RANDOM}};
  cache_41_5 = _RAND_415[15:0];
  _RAND_416 = {1{`RANDOM}};
  cache_41_6 = _RAND_416[15:0];
  _RAND_417 = {1{`RANDOM}};
  cache_41_7 = _RAND_417[15:0];
  _RAND_418 = {1{`RANDOM}};
  cache_41_8 = _RAND_418[15:0];
  _RAND_419 = {1{`RANDOM}};
  cache_41_9 = _RAND_419[15:0];
  _RAND_420 = {1{`RANDOM}};
  cache_42_0 = _RAND_420[15:0];
  _RAND_421 = {1{`RANDOM}};
  cache_42_1 = _RAND_421[15:0];
  _RAND_422 = {1{`RANDOM}};
  cache_42_2 = _RAND_422[15:0];
  _RAND_423 = {1{`RANDOM}};
  cache_42_3 = _RAND_423[15:0];
  _RAND_424 = {1{`RANDOM}};
  cache_42_4 = _RAND_424[15:0];
  _RAND_425 = {1{`RANDOM}};
  cache_42_5 = _RAND_425[15:0];
  _RAND_426 = {1{`RANDOM}};
  cache_42_6 = _RAND_426[15:0];
  _RAND_427 = {1{`RANDOM}};
  cache_42_7 = _RAND_427[15:0];
  _RAND_428 = {1{`RANDOM}};
  cache_42_8 = _RAND_428[15:0];
  _RAND_429 = {1{`RANDOM}};
  cache_42_9 = _RAND_429[15:0];
  _RAND_430 = {1{`RANDOM}};
  cache_43_0 = _RAND_430[15:0];
  _RAND_431 = {1{`RANDOM}};
  cache_43_1 = _RAND_431[15:0];
  _RAND_432 = {1{`RANDOM}};
  cache_43_2 = _RAND_432[15:0];
  _RAND_433 = {1{`RANDOM}};
  cache_43_3 = _RAND_433[15:0];
  _RAND_434 = {1{`RANDOM}};
  cache_43_4 = _RAND_434[15:0];
  _RAND_435 = {1{`RANDOM}};
  cache_43_5 = _RAND_435[15:0];
  _RAND_436 = {1{`RANDOM}};
  cache_43_6 = _RAND_436[15:0];
  _RAND_437 = {1{`RANDOM}};
  cache_43_7 = _RAND_437[15:0];
  _RAND_438 = {1{`RANDOM}};
  cache_43_8 = _RAND_438[15:0];
  _RAND_439 = {1{`RANDOM}};
  cache_43_9 = _RAND_439[15:0];
  _RAND_440 = {1{`RANDOM}};
  cache_44_0 = _RAND_440[15:0];
  _RAND_441 = {1{`RANDOM}};
  cache_44_1 = _RAND_441[15:0];
  _RAND_442 = {1{`RANDOM}};
  cache_44_2 = _RAND_442[15:0];
  _RAND_443 = {1{`RANDOM}};
  cache_44_3 = _RAND_443[15:0];
  _RAND_444 = {1{`RANDOM}};
  cache_44_4 = _RAND_444[15:0];
  _RAND_445 = {1{`RANDOM}};
  cache_44_5 = _RAND_445[15:0];
  _RAND_446 = {1{`RANDOM}};
  cache_44_6 = _RAND_446[15:0];
  _RAND_447 = {1{`RANDOM}};
  cache_44_7 = _RAND_447[15:0];
  _RAND_448 = {1{`RANDOM}};
  cache_44_8 = _RAND_448[15:0];
  _RAND_449 = {1{`RANDOM}};
  cache_44_9 = _RAND_449[15:0];
  _RAND_450 = {1{`RANDOM}};
  cache_45_0 = _RAND_450[15:0];
  _RAND_451 = {1{`RANDOM}};
  cache_45_1 = _RAND_451[15:0];
  _RAND_452 = {1{`RANDOM}};
  cache_45_2 = _RAND_452[15:0];
  _RAND_453 = {1{`RANDOM}};
  cache_45_3 = _RAND_453[15:0];
  _RAND_454 = {1{`RANDOM}};
  cache_45_4 = _RAND_454[15:0];
  _RAND_455 = {1{`RANDOM}};
  cache_45_5 = _RAND_455[15:0];
  _RAND_456 = {1{`RANDOM}};
  cache_45_6 = _RAND_456[15:0];
  _RAND_457 = {1{`RANDOM}};
  cache_45_7 = _RAND_457[15:0];
  _RAND_458 = {1{`RANDOM}};
  cache_45_8 = _RAND_458[15:0];
  _RAND_459 = {1{`RANDOM}};
  cache_45_9 = _RAND_459[15:0];
  _RAND_460 = {1{`RANDOM}};
  cache_46_0 = _RAND_460[15:0];
  _RAND_461 = {1{`RANDOM}};
  cache_46_1 = _RAND_461[15:0];
  _RAND_462 = {1{`RANDOM}};
  cache_46_2 = _RAND_462[15:0];
  _RAND_463 = {1{`RANDOM}};
  cache_46_3 = _RAND_463[15:0];
  _RAND_464 = {1{`RANDOM}};
  cache_46_4 = _RAND_464[15:0];
  _RAND_465 = {1{`RANDOM}};
  cache_46_5 = _RAND_465[15:0];
  _RAND_466 = {1{`RANDOM}};
  cache_46_6 = _RAND_466[15:0];
  _RAND_467 = {1{`RANDOM}};
  cache_46_7 = _RAND_467[15:0];
  _RAND_468 = {1{`RANDOM}};
  cache_46_8 = _RAND_468[15:0];
  _RAND_469 = {1{`RANDOM}};
  cache_46_9 = _RAND_469[15:0];
  _RAND_470 = {1{`RANDOM}};
  cache_47_0 = _RAND_470[15:0];
  _RAND_471 = {1{`RANDOM}};
  cache_47_1 = _RAND_471[15:0];
  _RAND_472 = {1{`RANDOM}};
  cache_47_2 = _RAND_472[15:0];
  _RAND_473 = {1{`RANDOM}};
  cache_47_3 = _RAND_473[15:0];
  _RAND_474 = {1{`RANDOM}};
  cache_47_4 = _RAND_474[15:0];
  _RAND_475 = {1{`RANDOM}};
  cache_47_5 = _RAND_475[15:0];
  _RAND_476 = {1{`RANDOM}};
  cache_47_6 = _RAND_476[15:0];
  _RAND_477 = {1{`RANDOM}};
  cache_47_7 = _RAND_477[15:0];
  _RAND_478 = {1{`RANDOM}};
  cache_47_8 = _RAND_478[15:0];
  _RAND_479 = {1{`RANDOM}};
  cache_47_9 = _RAND_479[15:0];
  _RAND_480 = {1{`RANDOM}};
  cache_48_0 = _RAND_480[15:0];
  _RAND_481 = {1{`RANDOM}};
  cache_48_1 = _RAND_481[15:0];
  _RAND_482 = {1{`RANDOM}};
  cache_48_2 = _RAND_482[15:0];
  _RAND_483 = {1{`RANDOM}};
  cache_48_3 = _RAND_483[15:0];
  _RAND_484 = {1{`RANDOM}};
  cache_48_4 = _RAND_484[15:0];
  _RAND_485 = {1{`RANDOM}};
  cache_48_5 = _RAND_485[15:0];
  _RAND_486 = {1{`RANDOM}};
  cache_48_6 = _RAND_486[15:0];
  _RAND_487 = {1{`RANDOM}};
  cache_48_7 = _RAND_487[15:0];
  _RAND_488 = {1{`RANDOM}};
  cache_48_8 = _RAND_488[15:0];
  _RAND_489 = {1{`RANDOM}};
  cache_48_9 = _RAND_489[15:0];
  _RAND_490 = {1{`RANDOM}};
  cache_49_0 = _RAND_490[15:0];
  _RAND_491 = {1{`RANDOM}};
  cache_49_1 = _RAND_491[15:0];
  _RAND_492 = {1{`RANDOM}};
  cache_49_2 = _RAND_492[15:0];
  _RAND_493 = {1{`RANDOM}};
  cache_49_3 = _RAND_493[15:0];
  _RAND_494 = {1{`RANDOM}};
  cache_49_4 = _RAND_494[15:0];
  _RAND_495 = {1{`RANDOM}};
  cache_49_5 = _RAND_495[15:0];
  _RAND_496 = {1{`RANDOM}};
  cache_49_6 = _RAND_496[15:0];
  _RAND_497 = {1{`RANDOM}};
  cache_49_7 = _RAND_497[15:0];
  _RAND_498 = {1{`RANDOM}};
  cache_49_8 = _RAND_498[15:0];
  _RAND_499 = {1{`RANDOM}};
  cache_49_9 = _RAND_499[15:0];
  _RAND_500 = {1{`RANDOM}};
  cache_50_0 = _RAND_500[15:0];
  _RAND_501 = {1{`RANDOM}};
  cache_50_1 = _RAND_501[15:0];
  _RAND_502 = {1{`RANDOM}};
  cache_50_2 = _RAND_502[15:0];
  _RAND_503 = {1{`RANDOM}};
  cache_50_3 = _RAND_503[15:0];
  _RAND_504 = {1{`RANDOM}};
  cache_50_4 = _RAND_504[15:0];
  _RAND_505 = {1{`RANDOM}};
  cache_50_5 = _RAND_505[15:0];
  _RAND_506 = {1{`RANDOM}};
  cache_50_6 = _RAND_506[15:0];
  _RAND_507 = {1{`RANDOM}};
  cache_50_7 = _RAND_507[15:0];
  _RAND_508 = {1{`RANDOM}};
  cache_50_8 = _RAND_508[15:0];
  _RAND_509 = {1{`RANDOM}};
  cache_50_9 = _RAND_509[15:0];
  _RAND_510 = {1{`RANDOM}};
  cache_51_0 = _RAND_510[15:0];
  _RAND_511 = {1{`RANDOM}};
  cache_51_1 = _RAND_511[15:0];
  _RAND_512 = {1{`RANDOM}};
  cache_51_2 = _RAND_512[15:0];
  _RAND_513 = {1{`RANDOM}};
  cache_51_3 = _RAND_513[15:0];
  _RAND_514 = {1{`RANDOM}};
  cache_51_4 = _RAND_514[15:0];
  _RAND_515 = {1{`RANDOM}};
  cache_51_5 = _RAND_515[15:0];
  _RAND_516 = {1{`RANDOM}};
  cache_51_6 = _RAND_516[15:0];
  _RAND_517 = {1{`RANDOM}};
  cache_51_7 = _RAND_517[15:0];
  _RAND_518 = {1{`RANDOM}};
  cache_51_8 = _RAND_518[15:0];
  _RAND_519 = {1{`RANDOM}};
  cache_51_9 = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  cache_52_0 = _RAND_520[15:0];
  _RAND_521 = {1{`RANDOM}};
  cache_52_1 = _RAND_521[15:0];
  _RAND_522 = {1{`RANDOM}};
  cache_52_2 = _RAND_522[15:0];
  _RAND_523 = {1{`RANDOM}};
  cache_52_3 = _RAND_523[15:0];
  _RAND_524 = {1{`RANDOM}};
  cache_52_4 = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  cache_52_5 = _RAND_525[15:0];
  _RAND_526 = {1{`RANDOM}};
  cache_52_6 = _RAND_526[15:0];
  _RAND_527 = {1{`RANDOM}};
  cache_52_7 = _RAND_527[15:0];
  _RAND_528 = {1{`RANDOM}};
  cache_52_8 = _RAND_528[15:0];
  _RAND_529 = {1{`RANDOM}};
  cache_52_9 = _RAND_529[15:0];
  _RAND_530 = {1{`RANDOM}};
  cache_53_0 = _RAND_530[15:0];
  _RAND_531 = {1{`RANDOM}};
  cache_53_1 = _RAND_531[15:0];
  _RAND_532 = {1{`RANDOM}};
  cache_53_2 = _RAND_532[15:0];
  _RAND_533 = {1{`RANDOM}};
  cache_53_3 = _RAND_533[15:0];
  _RAND_534 = {1{`RANDOM}};
  cache_53_4 = _RAND_534[15:0];
  _RAND_535 = {1{`RANDOM}};
  cache_53_5 = _RAND_535[15:0];
  _RAND_536 = {1{`RANDOM}};
  cache_53_6 = _RAND_536[15:0];
  _RAND_537 = {1{`RANDOM}};
  cache_53_7 = _RAND_537[15:0];
  _RAND_538 = {1{`RANDOM}};
  cache_53_8 = _RAND_538[15:0];
  _RAND_539 = {1{`RANDOM}};
  cache_53_9 = _RAND_539[15:0];
  _RAND_540 = {1{`RANDOM}};
  cache_54_0 = _RAND_540[15:0];
  _RAND_541 = {1{`RANDOM}};
  cache_54_1 = _RAND_541[15:0];
  _RAND_542 = {1{`RANDOM}};
  cache_54_2 = _RAND_542[15:0];
  _RAND_543 = {1{`RANDOM}};
  cache_54_3 = _RAND_543[15:0];
  _RAND_544 = {1{`RANDOM}};
  cache_54_4 = _RAND_544[15:0];
  _RAND_545 = {1{`RANDOM}};
  cache_54_5 = _RAND_545[15:0];
  _RAND_546 = {1{`RANDOM}};
  cache_54_6 = _RAND_546[15:0];
  _RAND_547 = {1{`RANDOM}};
  cache_54_7 = _RAND_547[15:0];
  _RAND_548 = {1{`RANDOM}};
  cache_54_8 = _RAND_548[15:0];
  _RAND_549 = {1{`RANDOM}};
  cache_54_9 = _RAND_549[15:0];
  _RAND_550 = {1{`RANDOM}};
  cache_55_0 = _RAND_550[15:0];
  _RAND_551 = {1{`RANDOM}};
  cache_55_1 = _RAND_551[15:0];
  _RAND_552 = {1{`RANDOM}};
  cache_55_2 = _RAND_552[15:0];
  _RAND_553 = {1{`RANDOM}};
  cache_55_3 = _RAND_553[15:0];
  _RAND_554 = {1{`RANDOM}};
  cache_55_4 = _RAND_554[15:0];
  _RAND_555 = {1{`RANDOM}};
  cache_55_5 = _RAND_555[15:0];
  _RAND_556 = {1{`RANDOM}};
  cache_55_6 = _RAND_556[15:0];
  _RAND_557 = {1{`RANDOM}};
  cache_55_7 = _RAND_557[15:0];
  _RAND_558 = {1{`RANDOM}};
  cache_55_8 = _RAND_558[15:0];
  _RAND_559 = {1{`RANDOM}};
  cache_55_9 = _RAND_559[15:0];
  _RAND_560 = {1{`RANDOM}};
  cache_56_0 = _RAND_560[15:0];
  _RAND_561 = {1{`RANDOM}};
  cache_56_1 = _RAND_561[15:0];
  _RAND_562 = {1{`RANDOM}};
  cache_56_2 = _RAND_562[15:0];
  _RAND_563 = {1{`RANDOM}};
  cache_56_3 = _RAND_563[15:0];
  _RAND_564 = {1{`RANDOM}};
  cache_56_4 = _RAND_564[15:0];
  _RAND_565 = {1{`RANDOM}};
  cache_56_5 = _RAND_565[15:0];
  _RAND_566 = {1{`RANDOM}};
  cache_56_6 = _RAND_566[15:0];
  _RAND_567 = {1{`RANDOM}};
  cache_56_7 = _RAND_567[15:0];
  _RAND_568 = {1{`RANDOM}};
  cache_56_8 = _RAND_568[15:0];
  _RAND_569 = {1{`RANDOM}};
  cache_56_9 = _RAND_569[15:0];
  _RAND_570 = {1{`RANDOM}};
  cache_57_0 = _RAND_570[15:0];
  _RAND_571 = {1{`RANDOM}};
  cache_57_1 = _RAND_571[15:0];
  _RAND_572 = {1{`RANDOM}};
  cache_57_2 = _RAND_572[15:0];
  _RAND_573 = {1{`RANDOM}};
  cache_57_3 = _RAND_573[15:0];
  _RAND_574 = {1{`RANDOM}};
  cache_57_4 = _RAND_574[15:0];
  _RAND_575 = {1{`RANDOM}};
  cache_57_5 = _RAND_575[15:0];
  _RAND_576 = {1{`RANDOM}};
  cache_57_6 = _RAND_576[15:0];
  _RAND_577 = {1{`RANDOM}};
  cache_57_7 = _RAND_577[15:0];
  _RAND_578 = {1{`RANDOM}};
  cache_57_8 = _RAND_578[15:0];
  _RAND_579 = {1{`RANDOM}};
  cache_57_9 = _RAND_579[15:0];
  _RAND_580 = {1{`RANDOM}};
  cache_58_0 = _RAND_580[15:0];
  _RAND_581 = {1{`RANDOM}};
  cache_58_1 = _RAND_581[15:0];
  _RAND_582 = {1{`RANDOM}};
  cache_58_2 = _RAND_582[15:0];
  _RAND_583 = {1{`RANDOM}};
  cache_58_3 = _RAND_583[15:0];
  _RAND_584 = {1{`RANDOM}};
  cache_58_4 = _RAND_584[15:0];
  _RAND_585 = {1{`RANDOM}};
  cache_58_5 = _RAND_585[15:0];
  _RAND_586 = {1{`RANDOM}};
  cache_58_6 = _RAND_586[15:0];
  _RAND_587 = {1{`RANDOM}};
  cache_58_7 = _RAND_587[15:0];
  _RAND_588 = {1{`RANDOM}};
  cache_58_8 = _RAND_588[15:0];
  _RAND_589 = {1{`RANDOM}};
  cache_58_9 = _RAND_589[15:0];
  _RAND_590 = {1{`RANDOM}};
  cache_59_0 = _RAND_590[15:0];
  _RAND_591 = {1{`RANDOM}};
  cache_59_1 = _RAND_591[15:0];
  _RAND_592 = {1{`RANDOM}};
  cache_59_2 = _RAND_592[15:0];
  _RAND_593 = {1{`RANDOM}};
  cache_59_3 = _RAND_593[15:0];
  _RAND_594 = {1{`RANDOM}};
  cache_59_4 = _RAND_594[15:0];
  _RAND_595 = {1{`RANDOM}};
  cache_59_5 = _RAND_595[15:0];
  _RAND_596 = {1{`RANDOM}};
  cache_59_6 = _RAND_596[15:0];
  _RAND_597 = {1{`RANDOM}};
  cache_59_7 = _RAND_597[15:0];
  _RAND_598 = {1{`RANDOM}};
  cache_59_8 = _RAND_598[15:0];
  _RAND_599 = {1{`RANDOM}};
  cache_59_9 = _RAND_599[15:0];
  _RAND_600 = {1{`RANDOM}};
  cache_60_0 = _RAND_600[15:0];
  _RAND_601 = {1{`RANDOM}};
  cache_60_1 = _RAND_601[15:0];
  _RAND_602 = {1{`RANDOM}};
  cache_60_2 = _RAND_602[15:0];
  _RAND_603 = {1{`RANDOM}};
  cache_60_3 = _RAND_603[15:0];
  _RAND_604 = {1{`RANDOM}};
  cache_60_4 = _RAND_604[15:0];
  _RAND_605 = {1{`RANDOM}};
  cache_60_5 = _RAND_605[15:0];
  _RAND_606 = {1{`RANDOM}};
  cache_60_6 = _RAND_606[15:0];
  _RAND_607 = {1{`RANDOM}};
  cache_60_7 = _RAND_607[15:0];
  _RAND_608 = {1{`RANDOM}};
  cache_60_8 = _RAND_608[15:0];
  _RAND_609 = {1{`RANDOM}};
  cache_60_9 = _RAND_609[15:0];
  _RAND_610 = {1{`RANDOM}};
  cache_61_0 = _RAND_610[15:0];
  _RAND_611 = {1{`RANDOM}};
  cache_61_1 = _RAND_611[15:0];
  _RAND_612 = {1{`RANDOM}};
  cache_61_2 = _RAND_612[15:0];
  _RAND_613 = {1{`RANDOM}};
  cache_61_3 = _RAND_613[15:0];
  _RAND_614 = {1{`RANDOM}};
  cache_61_4 = _RAND_614[15:0];
  _RAND_615 = {1{`RANDOM}};
  cache_61_5 = _RAND_615[15:0];
  _RAND_616 = {1{`RANDOM}};
  cache_61_6 = _RAND_616[15:0];
  _RAND_617 = {1{`RANDOM}};
  cache_61_7 = _RAND_617[15:0];
  _RAND_618 = {1{`RANDOM}};
  cache_61_8 = _RAND_618[15:0];
  _RAND_619 = {1{`RANDOM}};
  cache_61_9 = _RAND_619[15:0];
  _RAND_620 = {1{`RANDOM}};
  cache_62_0 = _RAND_620[15:0];
  _RAND_621 = {1{`RANDOM}};
  cache_62_1 = _RAND_621[15:0];
  _RAND_622 = {1{`RANDOM}};
  cache_62_2 = _RAND_622[15:0];
  _RAND_623 = {1{`RANDOM}};
  cache_62_3 = _RAND_623[15:0];
  _RAND_624 = {1{`RANDOM}};
  cache_62_4 = _RAND_624[15:0];
  _RAND_625 = {1{`RANDOM}};
  cache_62_5 = _RAND_625[15:0];
  _RAND_626 = {1{`RANDOM}};
  cache_62_6 = _RAND_626[15:0];
  _RAND_627 = {1{`RANDOM}};
  cache_62_7 = _RAND_627[15:0];
  _RAND_628 = {1{`RANDOM}};
  cache_62_8 = _RAND_628[15:0];
  _RAND_629 = {1{`RANDOM}};
  cache_62_9 = _RAND_629[15:0];
  _RAND_630 = {1{`RANDOM}};
  cache_63_0 = _RAND_630[15:0];
  _RAND_631 = {1{`RANDOM}};
  cache_63_1 = _RAND_631[15:0];
  _RAND_632 = {1{`RANDOM}};
  cache_63_2 = _RAND_632[15:0];
  _RAND_633 = {1{`RANDOM}};
  cache_63_3 = _RAND_633[15:0];
  _RAND_634 = {1{`RANDOM}};
  cache_63_4 = _RAND_634[15:0];
  _RAND_635 = {1{`RANDOM}};
  cache_63_5 = _RAND_635[15:0];
  _RAND_636 = {1{`RANDOM}};
  cache_63_6 = _RAND_636[15:0];
  _RAND_637 = {1{`RANDOM}};
  cache_63_7 = _RAND_637[15:0];
  _RAND_638 = {1{`RANDOM}};
  cache_63_8 = _RAND_638[15:0];
  _RAND_639 = {1{`RANDOM}};
  cache_63_9 = _RAND_639[15:0];
  _RAND_640 = {1{`RANDOM}};
  cnt_ic_ccnt = _RAND_640[9:0];
  _RAND_641 = {1{`RANDOM}};
  cnt_ic_cend = _RAND_641[9:0];
  _RAND_642 = {1{`RANDOM}};
  cnt_x_ccnt = _RAND_642[9:0];
  _RAND_643 = {1{`RANDOM}};
  cnt_x_cend = _RAND_643[9:0];
  _RAND_644 = {1{`RANDOM}};
  cnt_y_ccnt = _RAND_644[9:0];
  _RAND_645 = {1{`RANDOM}};
  cnt_y_cend = _RAND_645[9:0];
  _RAND_646 = {1{`RANDOM}};
  state = _RAND_646[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadSwitch(
  input         clock,
  input         reset,
  input         io_flag_job,
  input  [1:0]  io_job,
  input         io_valid_in,
  output        io_valid_out_calc8x8,
  input  [15:0] io_from_mat_0,
  input  [15:0] io_from_mat_1,
  input  [15:0] io_from_mat_2,
  input  [15:0] io_from_mat_3,
  input  [15:0] io_from_mat_4,
  input  [15:0] io_from_mat_5,
  input  [15:0] io_from_mat_6,
  input  [15:0] io_from_mat_7,
  input  [15:0] io_from_mat_8,
  input  [15:0] io_from_mat_9,
  input  [15:0] io_from_mat_10,
  input  [15:0] io_from_mat_11,
  input  [15:0] io_from_mat_12,
  input  [15:0] io_from_mat_13,
  input  [15:0] io_from_mat_14,
  input  [15:0] io_from_mat_15,
  input  [15:0] io_from_mat_16,
  input  [15:0] io_from_mat_17,
  input  [15:0] io_from_mat_18,
  input  [15:0] io_from_mat_19,
  input  [15:0] io_from_mat_20,
  input  [15:0] io_from_mat_21,
  input  [15:0] io_from_mat_22,
  input  [15:0] io_from_mat_23,
  input  [15:0] io_from_mat_24,
  input  [15:0] io_from_mat_25,
  input  [15:0] io_from_mat_26,
  input  [15:0] io_from_mat_27,
  input  [15:0] io_from_mat_28,
  input  [15:0] io_from_mat_29,
  input  [15:0] io_from_mat_30,
  input  [15:0] io_from_mat_31,
  input  [15:0] io_from_mat_32,
  input  [15:0] io_from_mat_33,
  input  [15:0] io_from_mat_34,
  input  [15:0] io_from_mat_35,
  input  [15:0] io_from_mat_36,
  input  [15:0] io_from_mat_37,
  input  [15:0] io_from_mat_38,
  input  [15:0] io_from_mat_39,
  input  [15:0] io_from_mat_40,
  input  [15:0] io_from_mat_41,
  input  [15:0] io_from_mat_42,
  input  [15:0] io_from_mat_43,
  input  [15:0] io_from_mat_44,
  input  [15:0] io_from_mat_45,
  input  [15:0] io_from_mat_46,
  input  [15:0] io_from_mat_47,
  input  [15:0] io_from_mat_48,
  input  [15:0] io_from_mat_49,
  input  [15:0] io_from_mat_50,
  input  [15:0] io_from_mat_51,
  input  [15:0] io_from_mat_52,
  input  [15:0] io_from_mat_53,
  input  [15:0] io_from_mat_54,
  input  [15:0] io_from_mat_55,
  input  [15:0] io_from_mat_56,
  input  [15:0] io_from_mat_57,
  input  [15:0] io_from_mat_58,
  input  [15:0] io_from_mat_59,
  input  [15:0] io_from_mat_60,
  input  [15:0] io_from_mat_61,
  input  [15:0] io_from_mat_62,
  input  [15:0] io_from_mat_63,
  input  [15:0] io_from_up_0,
  input  [15:0] io_from_up_1,
  input  [15:0] io_from_up_2,
  input  [15:0] io_from_up_3,
  input  [15:0] io_from_up_4,
  input  [15:0] io_from_up_5,
  input  [15:0] io_from_up_6,
  input  [15:0] io_from_up_7,
  input  [15:0] io_from_up_8,
  input  [15:0] io_from_up_9,
  input  [15:0] io_from_down_0,
  input  [15:0] io_from_down_1,
  input  [15:0] io_from_down_2,
  input  [15:0] io_from_down_3,
  input  [15:0] io_from_down_4,
  input  [15:0] io_from_down_5,
  input  [15:0] io_from_down_6,
  input  [15:0] io_from_down_7,
  input  [15:0] io_from_down_8,
  input  [15:0] io_from_down_9,
  input  [15:0] io_from_left_0,
  input  [15:0] io_from_left_1,
  input  [15:0] io_from_left_2,
  input  [15:0] io_from_left_3,
  input  [15:0] io_from_left_4,
  input  [15:0] io_from_left_5,
  input  [15:0] io_from_left_6,
  input  [15:0] io_from_left_7,
  input  [15:0] io_from_right_0,
  input  [15:0] io_from_right_1,
  input  [15:0] io_from_right_2,
  input  [15:0] io_from_right_3,
  input  [15:0] io_from_right_4,
  input  [15:0] io_from_right_5,
  input  [15:0] io_from_right_6,
  input  [15:0] io_from_right_7,
  input  [15:0] io_from_weight_0,
  input  [15:0] io_from_weight_1,
  input  [15:0] io_from_weight_2,
  input  [15:0] io_from_weight_3,
  input  [15:0] io_from_weight_4,
  input  [15:0] io_from_weight_5,
  input  [15:0] io_from_weight_6,
  input  [15:0] io_from_weight_7,
  input  [15:0] io_from_weight_8,
  output [15:0] io_to_calc8x8_mat_0,
  output [15:0] io_to_calc8x8_mat_1,
  output [15:0] io_to_calc8x8_mat_2,
  output [15:0] io_to_calc8x8_mat_3,
  output [15:0] io_to_calc8x8_mat_4,
  output [15:0] io_to_calc8x8_mat_5,
  output [15:0] io_to_calc8x8_mat_6,
  output [15:0] io_to_calc8x8_mat_7,
  output [15:0] io_to_calc8x8_mat_8,
  output [15:0] io_to_calc8x8_mat_9,
  output [15:0] io_to_calc8x8_mat_10,
  output [15:0] io_to_calc8x8_mat_11,
  output [15:0] io_to_calc8x8_mat_12,
  output [15:0] io_to_calc8x8_mat_13,
  output [15:0] io_to_calc8x8_mat_14,
  output [15:0] io_to_calc8x8_mat_15,
  output [15:0] io_to_calc8x8_mat_16,
  output [15:0] io_to_calc8x8_mat_17,
  output [15:0] io_to_calc8x8_mat_18,
  output [15:0] io_to_calc8x8_mat_19,
  output [15:0] io_to_calc8x8_mat_20,
  output [15:0] io_to_calc8x8_mat_21,
  output [15:0] io_to_calc8x8_mat_22,
  output [15:0] io_to_calc8x8_mat_23,
  output [15:0] io_to_calc8x8_mat_24,
  output [15:0] io_to_calc8x8_mat_25,
  output [15:0] io_to_calc8x8_mat_26,
  output [15:0] io_to_calc8x8_mat_27,
  output [15:0] io_to_calc8x8_mat_28,
  output [15:0] io_to_calc8x8_mat_29,
  output [15:0] io_to_calc8x8_mat_30,
  output [15:0] io_to_calc8x8_mat_31,
  output [15:0] io_to_calc8x8_mat_32,
  output [15:0] io_to_calc8x8_mat_33,
  output [15:0] io_to_calc8x8_mat_34,
  output [15:0] io_to_calc8x8_mat_35,
  output [15:0] io_to_calc8x8_mat_36,
  output [15:0] io_to_calc8x8_mat_37,
  output [15:0] io_to_calc8x8_mat_38,
  output [15:0] io_to_calc8x8_mat_39,
  output [15:0] io_to_calc8x8_mat_40,
  output [15:0] io_to_calc8x8_mat_41,
  output [15:0] io_to_calc8x8_mat_42,
  output [15:0] io_to_calc8x8_mat_43,
  output [15:0] io_to_calc8x8_mat_44,
  output [15:0] io_to_calc8x8_mat_45,
  output [15:0] io_to_calc8x8_mat_46,
  output [15:0] io_to_calc8x8_mat_47,
  output [15:0] io_to_calc8x8_mat_48,
  output [15:0] io_to_calc8x8_mat_49,
  output [15:0] io_to_calc8x8_mat_50,
  output [15:0] io_to_calc8x8_mat_51,
  output [15:0] io_to_calc8x8_mat_52,
  output [15:0] io_to_calc8x8_mat_53,
  output [15:0] io_to_calc8x8_mat_54,
  output [15:0] io_to_calc8x8_mat_55,
  output [15:0] io_to_calc8x8_mat_56,
  output [15:0] io_to_calc8x8_mat_57,
  output [15:0] io_to_calc8x8_mat_58,
  output [15:0] io_to_calc8x8_mat_59,
  output [15:0] io_to_calc8x8_mat_60,
  output [15:0] io_to_calc8x8_mat_61,
  output [15:0] io_to_calc8x8_mat_62,
  output [15:0] io_to_calc8x8_mat_63,
  output [15:0] io_to_calc8x8_up_0,
  output [15:0] io_to_calc8x8_up_1,
  output [15:0] io_to_calc8x8_up_2,
  output [15:0] io_to_calc8x8_up_3,
  output [15:0] io_to_calc8x8_up_4,
  output [15:0] io_to_calc8x8_up_5,
  output [15:0] io_to_calc8x8_up_6,
  output [15:0] io_to_calc8x8_up_7,
  output [15:0] io_to_calc8x8_up_8,
  output [15:0] io_to_calc8x8_up_9,
  output [15:0] io_to_calc8x8_down_0,
  output [15:0] io_to_calc8x8_down_1,
  output [15:0] io_to_calc8x8_down_2,
  output [15:0] io_to_calc8x8_down_3,
  output [15:0] io_to_calc8x8_down_4,
  output [15:0] io_to_calc8x8_down_5,
  output [15:0] io_to_calc8x8_down_6,
  output [15:0] io_to_calc8x8_down_7,
  output [15:0] io_to_calc8x8_down_8,
  output [15:0] io_to_calc8x8_down_9,
  output [15:0] io_to_calc8x8_left_0,
  output [15:0] io_to_calc8x8_left_1,
  output [15:0] io_to_calc8x8_left_2,
  output [15:0] io_to_calc8x8_left_3,
  output [15:0] io_to_calc8x8_left_4,
  output [15:0] io_to_calc8x8_left_5,
  output [15:0] io_to_calc8x8_left_6,
  output [15:0] io_to_calc8x8_left_7,
  output [15:0] io_to_calc8x8_right_0,
  output [15:0] io_to_calc8x8_right_1,
  output [15:0] io_to_calc8x8_right_2,
  output [15:0] io_to_calc8x8_right_3,
  output [15:0] io_to_calc8x8_right_4,
  output [15:0] io_to_calc8x8_right_5,
  output [15:0] io_to_calc8x8_right_6,
  output [15:0] io_to_calc8x8_right_7,
  output [15:0] io_to_weight_0_real_0,
  output [15:0] io_to_weight_0_real_1,
  output [15:0] io_to_weight_0_real_2,
  output [15:0] io_to_weight_0_real_3,
  output [15:0] io_to_weight_0_real_4,
  output [15:0] io_to_weight_0_real_5,
  output [15:0] io_to_weight_0_real_6,
  output [15:0] io_to_weight_0_real_7,
  output [15:0] io_to_weight_0_real_8,
  output [15:0] io_to_weight_0_real_9,
  output [15:0] io_to_weight_0_real_10,
  output [15:0] io_to_weight_0_real_11,
  output [15:0] io_to_weight_0_real_12,
  output [15:0] io_to_weight_0_real_13,
  output [15:0] io_to_weight_0_real_14,
  output [15:0] io_to_weight_0_real_15,
  output [15:0] io_to_weight_1_real_0,
  output [15:0] io_to_weight_1_real_1,
  output [15:0] io_to_weight_1_real_2,
  output [15:0] io_to_weight_1_real_3,
  output [15:0] io_to_weight_1_real_4,
  output [15:0] io_to_weight_1_real_5,
  output [15:0] io_to_weight_1_real_6,
  output [15:0] io_to_weight_1_real_7,
  output [15:0] io_to_weight_1_real_8,
  output [15:0] io_to_weight_1_real_9,
  output [15:0] io_to_weight_1_real_10,
  output [15:0] io_to_weight_1_real_11,
  output [15:0] io_to_weight_1_real_12,
  output [15:0] io_to_weight_1_real_13,
  output [15:0] io_to_weight_1_real_14,
  output [15:0] io_to_weight_1_real_15,
  output [15:0] io_to_weight_2_real_0,
  output [15:0] io_to_weight_2_real_1,
  output [15:0] io_to_weight_2_real_2,
  output [15:0] io_to_weight_2_real_3,
  output [15:0] io_to_weight_2_real_4,
  output [15:0] io_to_weight_2_real_5,
  output [15:0] io_to_weight_2_real_6,
  output [15:0] io_to_weight_2_real_7,
  output [15:0] io_to_weight_2_real_8,
  output [15:0] io_to_weight_2_real_9,
  output [15:0] io_to_weight_2_real_10,
  output [15:0] io_to_weight_2_real_11,
  output [15:0] io_to_weight_2_real_12,
  output [15:0] io_to_weight_2_real_13,
  output [15:0] io_to_weight_2_real_14,
  output [15:0] io_to_weight_2_real_15,
  output [15:0] io_to_weight_3_real_0,
  output [15:0] io_to_weight_3_real_1,
  output [15:0] io_to_weight_3_real_2,
  output [15:0] io_to_weight_3_real_3,
  output [15:0] io_to_weight_3_real_4,
  output [15:0] io_to_weight_3_real_5,
  output [15:0] io_to_weight_3_real_6,
  output [15:0] io_to_weight_3_real_7,
  output [15:0] io_to_weight_3_real_8,
  output [15:0] io_to_weight_3_real_9,
  output [15:0] io_to_weight_3_real_10,
  output [15:0] io_to_weight_3_real_11,
  output [15:0] io_to_weight_3_real_12,
  output [15:0] io_to_weight_3_real_13,
  output [15:0] io_to_weight_3_real_14,
  output [15:0] io_to_weight_3_real_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] job_type; // @[switch.scala 28:27]
  reg [15:0] cache_0; // @[switch.scala 30:24]
  reg [15:0] cache_1; // @[switch.scala 30:24]
  reg [15:0] cache_2; // @[switch.scala 30:24]
  reg [15:0] cache_3; // @[switch.scala 30:24]
  reg [15:0] cache_4; // @[switch.scala 30:24]
  reg [15:0] cache_5; // @[switch.scala 30:24]
  reg [15:0] cache_6; // @[switch.scala 30:24]
  reg [15:0] cache_7; // @[switch.scala 30:24]
  reg [15:0] cache_8; // @[switch.scala 30:24]
  reg [15:0] cache_9; // @[switch.scala 30:24]
  reg [15:0] cache_10; // @[switch.scala 30:24]
  reg [15:0] cache_11; // @[switch.scala 30:24]
  reg [15:0] cache_12; // @[switch.scala 30:24]
  reg [15:0] cache_13; // @[switch.scala 30:24]
  reg [15:0] cache_14; // @[switch.scala 30:24]
  reg [15:0] cache_15; // @[switch.scala 30:24]
  reg [15:0] cache_16; // @[switch.scala 30:24]
  reg [15:0] cache_17; // @[switch.scala 30:24]
  reg [15:0] cache_18; // @[switch.scala 30:24]
  reg [15:0] cache_19; // @[switch.scala 30:24]
  reg [15:0] cache_20; // @[switch.scala 30:24]
  reg [15:0] cache_21; // @[switch.scala 30:24]
  reg [15:0] cache_22; // @[switch.scala 30:24]
  reg [15:0] cache_23; // @[switch.scala 30:24]
  reg [15:0] cache_24; // @[switch.scala 30:24]
  reg [15:0] cache_25; // @[switch.scala 30:24]
  reg [15:0] cache_26; // @[switch.scala 30:24]
  reg [15:0] cache_27; // @[switch.scala 30:24]
  reg [15:0] cache_28; // @[switch.scala 30:24]
  reg [15:0] cache_29; // @[switch.scala 30:24]
  reg [15:0] cache_30; // @[switch.scala 30:24]
  reg [15:0] cache_31; // @[switch.scala 30:24]
  reg [15:0] cache_32; // @[switch.scala 30:24]
  reg [15:0] cache_33; // @[switch.scala 30:24]
  reg [15:0] cache_34; // @[switch.scala 30:24]
  reg [15:0] cache_35; // @[switch.scala 30:24]
  reg [15:0] cache_36; // @[switch.scala 30:24]
  reg [15:0] cache_37; // @[switch.scala 30:24]
  reg [15:0] cache_38; // @[switch.scala 30:24]
  reg [15:0] cache_39; // @[switch.scala 30:24]
  reg [15:0] cache_40; // @[switch.scala 30:24]
  reg [15:0] cache_41; // @[switch.scala 30:24]
  reg [15:0] cache_42; // @[switch.scala 30:24]
  reg [15:0] cache_43; // @[switch.scala 30:24]
  reg [15:0] cache_44; // @[switch.scala 30:24]
  reg [15:0] cache_45; // @[switch.scala 30:24]
  reg [15:0] cache_46; // @[switch.scala 30:24]
  reg [15:0] cache_47; // @[switch.scala 30:24]
  reg [15:0] cache_48; // @[switch.scala 30:24]
  reg [15:0] cache_49; // @[switch.scala 30:24]
  reg [15:0] cache_50; // @[switch.scala 30:24]
  reg [15:0] cache_51; // @[switch.scala 30:24]
  reg [15:0] cache_52; // @[switch.scala 30:24]
  reg [15:0] cache_53; // @[switch.scala 30:24]
  reg [15:0] cache_54; // @[switch.scala 30:24]
  reg [15:0] cache_55; // @[switch.scala 30:24]
  reg [15:0] cache_56; // @[switch.scala 30:24]
  reg [15:0] cache_57; // @[switch.scala 30:24]
  reg [15:0] cache_58; // @[switch.scala 30:24]
  reg [15:0] cache_59; // @[switch.scala 30:24]
  reg [15:0] cache_60; // @[switch.scala 30:24]
  reg [15:0] cache_61; // @[switch.scala 30:24]
  reg [15:0] cache_62; // @[switch.scala 30:24]
  reg [15:0] cache_63; // @[switch.scala 30:24]
  reg  state_ccnt; // @[switch.scala 31:24]
  reg  state_cend; // @[switch.scala 31:24]
  wire  _T_66 = 2'h1 == job_type; // @[Conditional.scala 37:30]
  wire  _T_69 = 2'h0 == job_type; // @[Conditional.scala 37:30]
  wire  _T_72 = 2'h2 == job_type; // @[Conditional.scala 37:30]
  wire  nxt = state_ccnt == state_cend; // @[utils.scala 17:20]
  wire  _state_ccnt_T_2 = nxt ? 1'h0 : state_ccnt + 1'h1; // @[utils.scala 18:20]
  wire [15:0] _GEN_1 = nxt ? $signed(io_from_right_0) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_2 = nxt ? $signed(io_from_right_1) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_3 = nxt ? $signed(io_from_right_2) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_4 = nxt ? $signed(io_from_right_3) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_5 = nxt ? $signed(io_from_right_4) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_6 = nxt ? $signed(io_from_right_5) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_7 = nxt ? $signed(io_from_right_6) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_8 = nxt ? $signed(io_from_right_7) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_9 = nxt ? $signed(io_from_left_0) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_10 = nxt ? $signed(io_from_left_1) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_11 = nxt ? $signed(io_from_left_2) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_12 = nxt ? $signed(io_from_left_3) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_13 = nxt ? $signed(io_from_left_4) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_14 = nxt ? $signed(io_from_left_5) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_15 = nxt ? $signed(io_from_left_6) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_16 = nxt ? $signed(io_from_left_7) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_17 = nxt ? $signed(io_from_down_0) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_18 = nxt ? $signed(io_from_down_1) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_19 = nxt ? $signed(io_from_down_2) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_20 = nxt ? $signed(io_from_down_3) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_21 = nxt ? $signed(io_from_down_4) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_22 = nxt ? $signed(io_from_down_5) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_23 = nxt ? $signed(io_from_down_6) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_24 = nxt ? $signed(io_from_down_7) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_25 = nxt ? $signed(io_from_down_8) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_26 = nxt ? $signed(io_from_down_9) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_27 = nxt ? $signed(io_from_up_0) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_28 = nxt ? $signed(io_from_up_1) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_29 = nxt ? $signed(io_from_up_2) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_30 = nxt ? $signed(io_from_up_3) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_31 = nxt ? $signed(io_from_up_4) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_32 = nxt ? $signed(io_from_up_5) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_33 = nxt ? $signed(io_from_up_6) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_34 = nxt ? $signed(io_from_up_7) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_35 = nxt ? $signed(io_from_up_8) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_36 = nxt ? $signed(io_from_up_9) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_37 = nxt ? $signed(io_from_mat_0) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_38 = nxt ? $signed(io_from_mat_1) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_39 = nxt ? $signed(io_from_mat_2) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_40 = nxt ? $signed(io_from_mat_3) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_41 = nxt ? $signed(io_from_mat_4) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_42 = nxt ? $signed(io_from_mat_5) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_43 = nxt ? $signed(io_from_mat_6) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_44 = nxt ? $signed(io_from_mat_7) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_45 = nxt ? $signed(io_from_mat_8) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_46 = nxt ? $signed(io_from_mat_9) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_47 = nxt ? $signed(io_from_mat_10) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_48 = nxt ? $signed(io_from_mat_11) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_49 = nxt ? $signed(io_from_mat_12) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_50 = nxt ? $signed(io_from_mat_13) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_51 = nxt ? $signed(io_from_mat_14) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_52 = nxt ? $signed(io_from_mat_15) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_53 = nxt ? $signed(io_from_mat_16) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_54 = nxt ? $signed(io_from_mat_17) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_55 = nxt ? $signed(io_from_mat_18) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_56 = nxt ? $signed(io_from_mat_19) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_57 = nxt ? $signed(io_from_mat_20) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_58 = nxt ? $signed(io_from_mat_21) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_59 = nxt ? $signed(io_from_mat_22) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_60 = nxt ? $signed(io_from_mat_23) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_61 = nxt ? $signed(io_from_mat_24) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_62 = nxt ? $signed(io_from_mat_25) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_63 = nxt ? $signed(io_from_mat_26) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_64 = nxt ? $signed(io_from_mat_27) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_65 = nxt ? $signed(io_from_mat_28) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_66 = nxt ? $signed(io_from_mat_29) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_67 = nxt ? $signed(io_from_mat_30) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_68 = nxt ? $signed(io_from_mat_31) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_69 = nxt ? $signed(io_from_mat_32) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_70 = nxt ? $signed(io_from_mat_33) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_71 = nxt ? $signed(io_from_mat_34) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_72 = nxt ? $signed(io_from_mat_35) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_73 = nxt ? $signed(io_from_mat_36) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_74 = nxt ? $signed(io_from_mat_37) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_75 = nxt ? $signed(io_from_mat_38) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_76 = nxt ? $signed(io_from_mat_39) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_77 = nxt ? $signed(io_from_mat_40) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_78 = nxt ? $signed(io_from_mat_41) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_79 = nxt ? $signed(io_from_mat_42) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_80 = nxt ? $signed(io_from_mat_43) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_81 = nxt ? $signed(io_from_mat_44) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_82 = nxt ? $signed(io_from_mat_45) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_83 = nxt ? $signed(io_from_mat_46) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_84 = nxt ? $signed(io_from_mat_47) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_85 = nxt ? $signed(io_from_mat_48) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_86 = nxt ? $signed(io_from_mat_49) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_87 = nxt ? $signed(io_from_mat_50) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_88 = nxt ? $signed(io_from_mat_51) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_89 = nxt ? $signed(io_from_mat_52) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_90 = nxt ? $signed(io_from_mat_53) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_91 = nxt ? $signed(io_from_mat_54) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_92 = nxt ? $signed(io_from_mat_55) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_93 = nxt ? $signed(io_from_mat_56) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_94 = nxt ? $signed(io_from_mat_57) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_95 = nxt ? $signed(io_from_mat_58) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_96 = nxt ? $signed(io_from_mat_59) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_97 = nxt ? $signed(io_from_mat_60) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_98 = nxt ? $signed(io_from_mat_61) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_99 = nxt ? $signed(io_from_mat_62) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_100 = nxt ? $signed(io_from_mat_63) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 57:35 switch.scala 35:19]
  wire [15:0] _GEN_101 = nxt ? $signed(cache_0) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_102 = nxt ? $signed(cache_1) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_103 = nxt ? $signed(cache_2) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_104 = nxt ? $signed(cache_3) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_105 = nxt ? $signed(cache_8) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_106 = nxt ? $signed(cache_9) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_107 = nxt ? $signed(cache_10) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_108 = nxt ? $signed(cache_11) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_109 = nxt ? $signed(cache_16) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_110 = nxt ? $signed(cache_17) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_111 = nxt ? $signed(cache_18) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_112 = nxt ? $signed(cache_19) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_113 = nxt ? $signed(cache_24) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_114 = nxt ? $signed(cache_25) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_115 = nxt ? $signed(cache_26) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_116 = nxt ? $signed(cache_27) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_117 = nxt ? $signed(cache_4) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_118 = nxt ? $signed(cache_5) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_119 = nxt ? $signed(cache_6) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_120 = nxt ? $signed(cache_7) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_121 = nxt ? $signed(cache_12) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_122 = nxt ? $signed(cache_13) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_123 = nxt ? $signed(cache_14) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_124 = nxt ? $signed(cache_15) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_125 = nxt ? $signed(cache_20) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_126 = nxt ? $signed(cache_21) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_127 = nxt ? $signed(cache_22) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_128 = nxt ? $signed(cache_23) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_129 = nxt ? $signed(cache_28) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_130 = nxt ? $signed(cache_29) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_131 = nxt ? $signed(cache_30) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_132 = nxt ? $signed(cache_31) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_133 = nxt ? $signed(cache_32) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_134 = nxt ? $signed(cache_33) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_135 = nxt ? $signed(cache_34) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_136 = nxt ? $signed(cache_35) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_137 = nxt ? $signed(cache_40) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_138 = nxt ? $signed(cache_41) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_139 = nxt ? $signed(cache_42) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_140 = nxt ? $signed(cache_43) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_141 = nxt ? $signed(cache_48) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_142 = nxt ? $signed(cache_49) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_143 = nxt ? $signed(cache_50) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_144 = nxt ? $signed(cache_51) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_145 = nxt ? $signed(cache_56) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_146 = nxt ? $signed(cache_57) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_147 = nxt ? $signed(cache_58) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_148 = nxt ? $signed(cache_59) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_149 = nxt ? $signed(cache_36) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_150 = nxt ? $signed(cache_37) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_151 = nxt ? $signed(cache_38) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_152 = nxt ? $signed(cache_39) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_153 = nxt ? $signed(cache_44) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_154 = nxt ? $signed(cache_45) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_155 = nxt ? $signed(cache_46) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_156 = nxt ? $signed(cache_47) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_157 = nxt ? $signed(cache_52) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_158 = nxt ? $signed(cache_53) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_159 = nxt ? $signed(cache_54) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_160 = nxt ? $signed(cache_55) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_161 = nxt ? $signed(cache_60) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_162 = nxt ? $signed(cache_61) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_163 = nxt ? $signed(cache_62) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_164 = nxt ? $signed(cache_63) : $signed(16'sh0); // @[switch.scala 55:34 switch.scala 62:71 switch.scala 36:18]
  wire [15:0] _GEN_165 = nxt ? $signed(cache_0) : $signed(io_from_mat_0); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_166 = nxt ? $signed(cache_1) : $signed(io_from_mat_1); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_167 = nxt ? $signed(cache_2) : $signed(io_from_mat_2); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_168 = nxt ? $signed(cache_3) : $signed(io_from_mat_3); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_169 = nxt ? $signed(cache_4) : $signed(io_from_mat_4); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_170 = nxt ? $signed(cache_5) : $signed(io_from_mat_5); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_171 = nxt ? $signed(cache_6) : $signed(io_from_mat_6); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_172 = nxt ? $signed(cache_7) : $signed(io_from_mat_7); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_173 = nxt ? $signed(cache_8) : $signed(io_from_mat_8); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_174 = nxt ? $signed(cache_9) : $signed(io_from_mat_9); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_175 = nxt ? $signed(cache_10) : $signed(io_from_mat_10); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_176 = nxt ? $signed(cache_11) : $signed(io_from_mat_11); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_177 = nxt ? $signed(cache_12) : $signed(io_from_mat_12); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_178 = nxt ? $signed(cache_13) : $signed(io_from_mat_13); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_179 = nxt ? $signed(cache_14) : $signed(io_from_mat_14); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_180 = nxt ? $signed(cache_15) : $signed(io_from_mat_15); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_181 = nxt ? $signed(cache_16) : $signed(io_from_mat_16); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_182 = nxt ? $signed(cache_17) : $signed(io_from_mat_17); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_183 = nxt ? $signed(cache_18) : $signed(io_from_mat_18); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_184 = nxt ? $signed(cache_19) : $signed(io_from_mat_19); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_185 = nxt ? $signed(cache_20) : $signed(io_from_mat_20); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_186 = nxt ? $signed(cache_21) : $signed(io_from_mat_21); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_187 = nxt ? $signed(cache_22) : $signed(io_from_mat_22); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_188 = nxt ? $signed(cache_23) : $signed(io_from_mat_23); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_189 = nxt ? $signed(cache_24) : $signed(io_from_mat_24); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_190 = nxt ? $signed(cache_25) : $signed(io_from_mat_25); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_191 = nxt ? $signed(cache_26) : $signed(io_from_mat_26); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_192 = nxt ? $signed(cache_27) : $signed(io_from_mat_27); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_193 = nxt ? $signed(cache_28) : $signed(io_from_mat_28); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_194 = nxt ? $signed(cache_29) : $signed(io_from_mat_29); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_195 = nxt ? $signed(cache_30) : $signed(io_from_mat_30); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_196 = nxt ? $signed(cache_31) : $signed(io_from_mat_31); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_197 = nxt ? $signed(cache_32) : $signed(io_from_mat_32); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_198 = nxt ? $signed(cache_33) : $signed(io_from_mat_33); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_199 = nxt ? $signed(cache_34) : $signed(io_from_mat_34); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_200 = nxt ? $signed(cache_35) : $signed(io_from_mat_35); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_201 = nxt ? $signed(cache_36) : $signed(io_from_mat_36); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_202 = nxt ? $signed(cache_37) : $signed(io_from_mat_37); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_203 = nxt ? $signed(cache_38) : $signed(io_from_mat_38); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_204 = nxt ? $signed(cache_39) : $signed(io_from_mat_39); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_205 = nxt ? $signed(cache_40) : $signed(io_from_mat_40); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_206 = nxt ? $signed(cache_41) : $signed(io_from_mat_41); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_207 = nxt ? $signed(cache_42) : $signed(io_from_mat_42); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_208 = nxt ? $signed(cache_43) : $signed(io_from_mat_43); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_209 = nxt ? $signed(cache_44) : $signed(io_from_mat_44); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_210 = nxt ? $signed(cache_45) : $signed(io_from_mat_45); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_211 = nxt ? $signed(cache_46) : $signed(io_from_mat_46); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_212 = nxt ? $signed(cache_47) : $signed(io_from_mat_47); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_213 = nxt ? $signed(cache_48) : $signed(io_from_mat_48); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_214 = nxt ? $signed(cache_49) : $signed(io_from_mat_49); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_215 = nxt ? $signed(cache_50) : $signed(io_from_mat_50); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_216 = nxt ? $signed(cache_51) : $signed(io_from_mat_51); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_217 = nxt ? $signed(cache_52) : $signed(io_from_mat_52); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_218 = nxt ? $signed(cache_53) : $signed(io_from_mat_53); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_219 = nxt ? $signed(cache_54) : $signed(io_from_mat_54); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_220 = nxt ? $signed(cache_55) : $signed(io_from_mat_55); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_221 = nxt ? $signed(cache_56) : $signed(io_from_mat_56); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_222 = nxt ? $signed(cache_57) : $signed(io_from_mat_57); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_223 = nxt ? $signed(cache_58) : $signed(io_from_mat_58); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_224 = nxt ? $signed(cache_59) : $signed(io_from_mat_59); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_225 = nxt ? $signed(cache_60) : $signed(io_from_mat_60); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_226 = nxt ? $signed(cache_61) : $signed(io_from_mat_61); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_227 = nxt ? $signed(cache_62) : $signed(io_from_mat_62); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire [15:0] _GEN_228 = nxt ? $signed(cache_63) : $signed(io_from_mat_63); // @[switch.scala 55:34 switch.scala 30:24 switch.scala 64:27]
  wire  _GEN_229 = _T_72 ? _state_ccnt_T_2 : state_ccnt; // @[Conditional.scala 39:67 utils.scala 18:14 switch.scala 31:24]
  wire [15:0] _GEN_231 = _T_72 ? $signed(_GEN_1) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_232 = _T_72 ? $signed(_GEN_2) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_233 = _T_72 ? $signed(_GEN_3) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_234 = _T_72 ? $signed(_GEN_4) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_235 = _T_72 ? $signed(_GEN_5) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_236 = _T_72 ? $signed(_GEN_6) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_237 = _T_72 ? $signed(_GEN_7) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_238 = _T_72 ? $signed(_GEN_8) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_239 = _T_72 ? $signed(_GEN_9) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_240 = _T_72 ? $signed(_GEN_10) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_241 = _T_72 ? $signed(_GEN_11) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_242 = _T_72 ? $signed(_GEN_12) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_243 = _T_72 ? $signed(_GEN_13) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_244 = _T_72 ? $signed(_GEN_14) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_245 = _T_72 ? $signed(_GEN_15) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_246 = _T_72 ? $signed(_GEN_16) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_247 = _T_72 ? $signed(_GEN_17) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_248 = _T_72 ? $signed(_GEN_18) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_249 = _T_72 ? $signed(_GEN_19) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_250 = _T_72 ? $signed(_GEN_20) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_251 = _T_72 ? $signed(_GEN_21) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_252 = _T_72 ? $signed(_GEN_22) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_253 = _T_72 ? $signed(_GEN_23) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_254 = _T_72 ? $signed(_GEN_24) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_255 = _T_72 ? $signed(_GEN_25) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_256 = _T_72 ? $signed(_GEN_26) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_257 = _T_72 ? $signed(_GEN_27) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_258 = _T_72 ? $signed(_GEN_28) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_259 = _T_72 ? $signed(_GEN_29) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_260 = _T_72 ? $signed(_GEN_30) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_261 = _T_72 ? $signed(_GEN_31) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_262 = _T_72 ? $signed(_GEN_32) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_263 = _T_72 ? $signed(_GEN_33) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_264 = _T_72 ? $signed(_GEN_34) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_265 = _T_72 ? $signed(_GEN_35) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_266 = _T_72 ? $signed(_GEN_36) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_267 = _T_72 ? $signed(_GEN_37) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_268 = _T_72 ? $signed(_GEN_38) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_269 = _T_72 ? $signed(_GEN_39) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_270 = _T_72 ? $signed(_GEN_40) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_271 = _T_72 ? $signed(_GEN_41) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_272 = _T_72 ? $signed(_GEN_42) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_273 = _T_72 ? $signed(_GEN_43) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_274 = _T_72 ? $signed(_GEN_44) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_275 = _T_72 ? $signed(_GEN_45) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_276 = _T_72 ? $signed(_GEN_46) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_277 = _T_72 ? $signed(_GEN_47) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_278 = _T_72 ? $signed(_GEN_48) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_279 = _T_72 ? $signed(_GEN_49) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_280 = _T_72 ? $signed(_GEN_50) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_281 = _T_72 ? $signed(_GEN_51) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_282 = _T_72 ? $signed(_GEN_52) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_283 = _T_72 ? $signed(_GEN_53) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_284 = _T_72 ? $signed(_GEN_54) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_285 = _T_72 ? $signed(_GEN_55) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_286 = _T_72 ? $signed(_GEN_56) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_287 = _T_72 ? $signed(_GEN_57) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_288 = _T_72 ? $signed(_GEN_58) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_289 = _T_72 ? $signed(_GEN_59) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_290 = _T_72 ? $signed(_GEN_60) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_291 = _T_72 ? $signed(_GEN_61) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_292 = _T_72 ? $signed(_GEN_62) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_293 = _T_72 ? $signed(_GEN_63) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_294 = _T_72 ? $signed(_GEN_64) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_295 = _T_72 ? $signed(_GEN_65) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_296 = _T_72 ? $signed(_GEN_66) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_297 = _T_72 ? $signed(_GEN_67) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_298 = _T_72 ? $signed(_GEN_68) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_299 = _T_72 ? $signed(_GEN_69) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_300 = _T_72 ? $signed(_GEN_70) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_301 = _T_72 ? $signed(_GEN_71) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_302 = _T_72 ? $signed(_GEN_72) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_303 = _T_72 ? $signed(_GEN_73) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_304 = _T_72 ? $signed(_GEN_74) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_305 = _T_72 ? $signed(_GEN_75) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_306 = _T_72 ? $signed(_GEN_76) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_307 = _T_72 ? $signed(_GEN_77) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_308 = _T_72 ? $signed(_GEN_78) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_309 = _T_72 ? $signed(_GEN_79) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_310 = _T_72 ? $signed(_GEN_80) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_311 = _T_72 ? $signed(_GEN_81) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_312 = _T_72 ? $signed(_GEN_82) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_313 = _T_72 ? $signed(_GEN_83) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_314 = _T_72 ? $signed(_GEN_84) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_315 = _T_72 ? $signed(_GEN_85) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_316 = _T_72 ? $signed(_GEN_86) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_317 = _T_72 ? $signed(_GEN_87) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_318 = _T_72 ? $signed(_GEN_88) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_319 = _T_72 ? $signed(_GEN_89) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_320 = _T_72 ? $signed(_GEN_90) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_321 = _T_72 ? $signed(_GEN_91) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_322 = _T_72 ? $signed(_GEN_92) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_323 = _T_72 ? $signed(_GEN_93) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_324 = _T_72 ? $signed(_GEN_94) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_325 = _T_72 ? $signed(_GEN_95) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_326 = _T_72 ? $signed(_GEN_96) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_327 = _T_72 ? $signed(_GEN_97) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_328 = _T_72 ? $signed(_GEN_98) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_329 = _T_72 ? $signed(_GEN_99) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_330 = _T_72 ? $signed(_GEN_100) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_331 = _T_72 ? $signed(_GEN_101) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_332 = _T_72 ? $signed(_GEN_102) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_333 = _T_72 ? $signed(_GEN_103) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_334 = _T_72 ? $signed(_GEN_104) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_335 = _T_72 ? $signed(_GEN_105) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_336 = _T_72 ? $signed(_GEN_106) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_337 = _T_72 ? $signed(_GEN_107) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_338 = _T_72 ? $signed(_GEN_108) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_339 = _T_72 ? $signed(_GEN_109) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_340 = _T_72 ? $signed(_GEN_110) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_341 = _T_72 ? $signed(_GEN_111) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_342 = _T_72 ? $signed(_GEN_112) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_343 = _T_72 ? $signed(_GEN_113) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_344 = _T_72 ? $signed(_GEN_114) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_345 = _T_72 ? $signed(_GEN_115) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_346 = _T_72 ? $signed(_GEN_116) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_347 = _T_72 ? $signed(_GEN_117) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_348 = _T_72 ? $signed(_GEN_118) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_349 = _T_72 ? $signed(_GEN_119) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_350 = _T_72 ? $signed(_GEN_120) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_351 = _T_72 ? $signed(_GEN_121) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_352 = _T_72 ? $signed(_GEN_122) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_353 = _T_72 ? $signed(_GEN_123) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_354 = _T_72 ? $signed(_GEN_124) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_355 = _T_72 ? $signed(_GEN_125) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_356 = _T_72 ? $signed(_GEN_126) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_357 = _T_72 ? $signed(_GEN_127) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_358 = _T_72 ? $signed(_GEN_128) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_359 = _T_72 ? $signed(_GEN_129) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_360 = _T_72 ? $signed(_GEN_130) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_361 = _T_72 ? $signed(_GEN_131) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_362 = _T_72 ? $signed(_GEN_132) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_363 = _T_72 ? $signed(_GEN_133) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_364 = _T_72 ? $signed(_GEN_134) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_365 = _T_72 ? $signed(_GEN_135) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_366 = _T_72 ? $signed(_GEN_136) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_367 = _T_72 ? $signed(_GEN_137) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_368 = _T_72 ? $signed(_GEN_138) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_369 = _T_72 ? $signed(_GEN_139) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_370 = _T_72 ? $signed(_GEN_140) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_371 = _T_72 ? $signed(_GEN_141) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_372 = _T_72 ? $signed(_GEN_142) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_373 = _T_72 ? $signed(_GEN_143) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_374 = _T_72 ? $signed(_GEN_144) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_375 = _T_72 ? $signed(_GEN_145) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_376 = _T_72 ? $signed(_GEN_146) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_377 = _T_72 ? $signed(_GEN_147) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_378 = _T_72 ? $signed(_GEN_148) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_379 = _T_72 ? $signed(_GEN_149) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_380 = _T_72 ? $signed(_GEN_150) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_381 = _T_72 ? $signed(_GEN_151) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_382 = _T_72 ? $signed(_GEN_152) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_383 = _T_72 ? $signed(_GEN_153) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_384 = _T_72 ? $signed(_GEN_154) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_385 = _T_72 ? $signed(_GEN_155) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_386 = _T_72 ? $signed(_GEN_156) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_387 = _T_72 ? $signed(_GEN_157) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_388 = _T_72 ? $signed(_GEN_158) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_389 = _T_72 ? $signed(_GEN_159) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_390 = _T_72 ? $signed(_GEN_160) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_391 = _T_72 ? $signed(_GEN_161) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_392 = _T_72 ? $signed(_GEN_162) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_393 = _T_72 ? $signed(_GEN_163) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_394 = _T_72 ? $signed(_GEN_164) : $signed(16'sh0); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_395 = _T_72 ? $signed(_GEN_165) : $signed(cache_0); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_396 = _T_72 ? $signed(_GEN_166) : $signed(cache_1); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_397 = _T_72 ? $signed(_GEN_167) : $signed(cache_2); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_398 = _T_72 ? $signed(_GEN_168) : $signed(cache_3); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_399 = _T_72 ? $signed(_GEN_169) : $signed(cache_4); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_400 = _T_72 ? $signed(_GEN_170) : $signed(cache_5); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_401 = _T_72 ? $signed(_GEN_171) : $signed(cache_6); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_402 = _T_72 ? $signed(_GEN_172) : $signed(cache_7); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_403 = _T_72 ? $signed(_GEN_173) : $signed(cache_8); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_404 = _T_72 ? $signed(_GEN_174) : $signed(cache_9); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_405 = _T_72 ? $signed(_GEN_175) : $signed(cache_10); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_406 = _T_72 ? $signed(_GEN_176) : $signed(cache_11); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_407 = _T_72 ? $signed(_GEN_177) : $signed(cache_12); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_408 = _T_72 ? $signed(_GEN_178) : $signed(cache_13); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_409 = _T_72 ? $signed(_GEN_179) : $signed(cache_14); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_410 = _T_72 ? $signed(_GEN_180) : $signed(cache_15); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_411 = _T_72 ? $signed(_GEN_181) : $signed(cache_16); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_412 = _T_72 ? $signed(_GEN_182) : $signed(cache_17); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_413 = _T_72 ? $signed(_GEN_183) : $signed(cache_18); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_414 = _T_72 ? $signed(_GEN_184) : $signed(cache_19); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_415 = _T_72 ? $signed(_GEN_185) : $signed(cache_20); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_416 = _T_72 ? $signed(_GEN_186) : $signed(cache_21); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_417 = _T_72 ? $signed(_GEN_187) : $signed(cache_22); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_418 = _T_72 ? $signed(_GEN_188) : $signed(cache_23); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_419 = _T_72 ? $signed(_GEN_189) : $signed(cache_24); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_420 = _T_72 ? $signed(_GEN_190) : $signed(cache_25); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_421 = _T_72 ? $signed(_GEN_191) : $signed(cache_26); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_422 = _T_72 ? $signed(_GEN_192) : $signed(cache_27); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_423 = _T_72 ? $signed(_GEN_193) : $signed(cache_28); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_424 = _T_72 ? $signed(_GEN_194) : $signed(cache_29); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_425 = _T_72 ? $signed(_GEN_195) : $signed(cache_30); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_426 = _T_72 ? $signed(_GEN_196) : $signed(cache_31); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_427 = _T_72 ? $signed(_GEN_197) : $signed(cache_32); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_428 = _T_72 ? $signed(_GEN_198) : $signed(cache_33); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_429 = _T_72 ? $signed(_GEN_199) : $signed(cache_34); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_430 = _T_72 ? $signed(_GEN_200) : $signed(cache_35); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_431 = _T_72 ? $signed(_GEN_201) : $signed(cache_36); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_432 = _T_72 ? $signed(_GEN_202) : $signed(cache_37); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_433 = _T_72 ? $signed(_GEN_203) : $signed(cache_38); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_434 = _T_72 ? $signed(_GEN_204) : $signed(cache_39); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_435 = _T_72 ? $signed(_GEN_205) : $signed(cache_40); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_436 = _T_72 ? $signed(_GEN_206) : $signed(cache_41); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_437 = _T_72 ? $signed(_GEN_207) : $signed(cache_42); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_438 = _T_72 ? $signed(_GEN_208) : $signed(cache_43); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_439 = _T_72 ? $signed(_GEN_209) : $signed(cache_44); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_440 = _T_72 ? $signed(_GEN_210) : $signed(cache_45); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_441 = _T_72 ? $signed(_GEN_211) : $signed(cache_46); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_442 = _T_72 ? $signed(_GEN_212) : $signed(cache_47); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_443 = _T_72 ? $signed(_GEN_213) : $signed(cache_48); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_444 = _T_72 ? $signed(_GEN_214) : $signed(cache_49); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_445 = _T_72 ? $signed(_GEN_215) : $signed(cache_50); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_446 = _T_72 ? $signed(_GEN_216) : $signed(cache_51); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_447 = _T_72 ? $signed(_GEN_217) : $signed(cache_52); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_448 = _T_72 ? $signed(_GEN_218) : $signed(cache_53); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_449 = _T_72 ? $signed(_GEN_219) : $signed(cache_54); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_450 = _T_72 ? $signed(_GEN_220) : $signed(cache_55); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_451 = _T_72 ? $signed(_GEN_221) : $signed(cache_56); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_452 = _T_72 ? $signed(_GEN_222) : $signed(cache_57); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_453 = _T_72 ? $signed(_GEN_223) : $signed(cache_58); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_454 = _T_72 ? $signed(_GEN_224) : $signed(cache_59); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_455 = _T_72 ? $signed(_GEN_225) : $signed(cache_60); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_456 = _T_72 ? $signed(_GEN_226) : $signed(cache_61); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_457 = _T_72 ? $signed(_GEN_227) : $signed(cache_62); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_458 = _T_72 ? $signed(_GEN_228) : $signed(cache_63); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire  _GEN_524 = _T_69 ? state_ccnt : _GEN_229; // @[Conditional.scala 39:67 switch.scala 31:24]
  wire  _GEN_525 = _T_69 ? 1'h0 : _T_72 & nxt; // @[Conditional.scala 39:67 switch.scala 33:26]
  wire [15:0] _GEN_526 = _T_69 ? $signed(16'sh0) : $signed(_GEN_231); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_527 = _T_69 ? $signed(16'sh0) : $signed(_GEN_232); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_528 = _T_69 ? $signed(16'sh0) : $signed(_GEN_233); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_529 = _T_69 ? $signed(16'sh0) : $signed(_GEN_234); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_530 = _T_69 ? $signed(16'sh0) : $signed(_GEN_235); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_531 = _T_69 ? $signed(16'sh0) : $signed(_GEN_236); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_532 = _T_69 ? $signed(16'sh0) : $signed(_GEN_237); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_533 = _T_69 ? $signed(16'sh0) : $signed(_GEN_238); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_534 = _T_69 ? $signed(16'sh0) : $signed(_GEN_239); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_535 = _T_69 ? $signed(16'sh0) : $signed(_GEN_240); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_536 = _T_69 ? $signed(16'sh0) : $signed(_GEN_241); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_537 = _T_69 ? $signed(16'sh0) : $signed(_GEN_242); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_538 = _T_69 ? $signed(16'sh0) : $signed(_GEN_243); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_539 = _T_69 ? $signed(16'sh0) : $signed(_GEN_244); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_540 = _T_69 ? $signed(16'sh0) : $signed(_GEN_245); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_541 = _T_69 ? $signed(16'sh0) : $signed(_GEN_246); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_542 = _T_69 ? $signed(16'sh0) : $signed(_GEN_247); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_543 = _T_69 ? $signed(16'sh0) : $signed(_GEN_248); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_544 = _T_69 ? $signed(16'sh0) : $signed(_GEN_249); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_545 = _T_69 ? $signed(16'sh0) : $signed(_GEN_250); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_546 = _T_69 ? $signed(16'sh0) : $signed(_GEN_251); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_547 = _T_69 ? $signed(16'sh0) : $signed(_GEN_252); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_548 = _T_69 ? $signed(16'sh0) : $signed(_GEN_253); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_549 = _T_69 ? $signed(16'sh0) : $signed(_GEN_254); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_550 = _T_69 ? $signed(16'sh0) : $signed(_GEN_255); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_551 = _T_69 ? $signed(16'sh0) : $signed(_GEN_256); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_552 = _T_69 ? $signed(16'sh0) : $signed(_GEN_257); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_553 = _T_69 ? $signed(16'sh0) : $signed(_GEN_258); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_554 = _T_69 ? $signed(16'sh0) : $signed(_GEN_259); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_555 = _T_69 ? $signed(16'sh0) : $signed(_GEN_260); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_556 = _T_69 ? $signed(16'sh0) : $signed(_GEN_261); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_557 = _T_69 ? $signed(16'sh0) : $signed(_GEN_262); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_558 = _T_69 ? $signed(16'sh0) : $signed(_GEN_263); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_559 = _T_69 ? $signed(16'sh0) : $signed(_GEN_264); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_560 = _T_69 ? $signed(16'sh0) : $signed(_GEN_265); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_561 = _T_69 ? $signed(16'sh0) : $signed(_GEN_266); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_562 = _T_69 ? $signed(16'sh0) : $signed(_GEN_267); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_563 = _T_69 ? $signed(16'sh0) : $signed(_GEN_268); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_564 = _T_69 ? $signed(16'sh0) : $signed(_GEN_269); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_565 = _T_69 ? $signed(16'sh0) : $signed(_GEN_270); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_566 = _T_69 ? $signed(16'sh0) : $signed(_GEN_271); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_567 = _T_69 ? $signed(16'sh0) : $signed(_GEN_272); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_568 = _T_69 ? $signed(16'sh0) : $signed(_GEN_273); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_569 = _T_69 ? $signed(16'sh0) : $signed(_GEN_274); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_570 = _T_69 ? $signed(16'sh0) : $signed(_GEN_275); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_571 = _T_69 ? $signed(16'sh0) : $signed(_GEN_276); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_572 = _T_69 ? $signed(16'sh0) : $signed(_GEN_277); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_573 = _T_69 ? $signed(16'sh0) : $signed(_GEN_278); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_574 = _T_69 ? $signed(16'sh0) : $signed(_GEN_279); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_575 = _T_69 ? $signed(16'sh0) : $signed(_GEN_280); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_576 = _T_69 ? $signed(16'sh0) : $signed(_GEN_281); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_577 = _T_69 ? $signed(16'sh0) : $signed(_GEN_282); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_578 = _T_69 ? $signed(16'sh0) : $signed(_GEN_283); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_579 = _T_69 ? $signed(16'sh0) : $signed(_GEN_284); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_580 = _T_69 ? $signed(16'sh0) : $signed(_GEN_285); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_581 = _T_69 ? $signed(16'sh0) : $signed(_GEN_286); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_582 = _T_69 ? $signed(16'sh0) : $signed(_GEN_287); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_583 = _T_69 ? $signed(16'sh0) : $signed(_GEN_288); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_584 = _T_69 ? $signed(16'sh0) : $signed(_GEN_289); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_585 = _T_69 ? $signed(16'sh0) : $signed(_GEN_290); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_586 = _T_69 ? $signed(16'sh0) : $signed(_GEN_291); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_587 = _T_69 ? $signed(16'sh0) : $signed(_GEN_292); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_588 = _T_69 ? $signed(16'sh0) : $signed(_GEN_293); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_589 = _T_69 ? $signed(16'sh0) : $signed(_GEN_294); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_590 = _T_69 ? $signed(16'sh0) : $signed(_GEN_295); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_591 = _T_69 ? $signed(16'sh0) : $signed(_GEN_296); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_592 = _T_69 ? $signed(16'sh0) : $signed(_GEN_297); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_593 = _T_69 ? $signed(16'sh0) : $signed(_GEN_298); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_594 = _T_69 ? $signed(16'sh0) : $signed(_GEN_299); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_595 = _T_69 ? $signed(16'sh0) : $signed(_GEN_300); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_596 = _T_69 ? $signed(16'sh0) : $signed(_GEN_301); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_597 = _T_69 ? $signed(16'sh0) : $signed(_GEN_302); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_598 = _T_69 ? $signed(16'sh0) : $signed(_GEN_303); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_599 = _T_69 ? $signed(16'sh0) : $signed(_GEN_304); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_600 = _T_69 ? $signed(16'sh0) : $signed(_GEN_305); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_601 = _T_69 ? $signed(16'sh0) : $signed(_GEN_306); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_602 = _T_69 ? $signed(16'sh0) : $signed(_GEN_307); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_603 = _T_69 ? $signed(16'sh0) : $signed(_GEN_308); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_604 = _T_69 ? $signed(16'sh0) : $signed(_GEN_309); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_605 = _T_69 ? $signed(16'sh0) : $signed(_GEN_310); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_606 = _T_69 ? $signed(16'sh0) : $signed(_GEN_311); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_607 = _T_69 ? $signed(16'sh0) : $signed(_GEN_312); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_608 = _T_69 ? $signed(16'sh0) : $signed(_GEN_313); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_609 = _T_69 ? $signed(16'sh0) : $signed(_GEN_314); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_610 = _T_69 ? $signed(16'sh0) : $signed(_GEN_315); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_611 = _T_69 ? $signed(16'sh0) : $signed(_GEN_316); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_612 = _T_69 ? $signed(16'sh0) : $signed(_GEN_317); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_613 = _T_69 ? $signed(16'sh0) : $signed(_GEN_318); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_614 = _T_69 ? $signed(16'sh0) : $signed(_GEN_319); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_615 = _T_69 ? $signed(16'sh0) : $signed(_GEN_320); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_616 = _T_69 ? $signed(16'sh0) : $signed(_GEN_321); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_617 = _T_69 ? $signed(16'sh0) : $signed(_GEN_322); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_618 = _T_69 ? $signed(16'sh0) : $signed(_GEN_323); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_619 = _T_69 ? $signed(16'sh0) : $signed(_GEN_324); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_620 = _T_69 ? $signed(16'sh0) : $signed(_GEN_325); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_621 = _T_69 ? $signed(16'sh0) : $signed(_GEN_326); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_622 = _T_69 ? $signed(16'sh0) : $signed(_GEN_327); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_623 = _T_69 ? $signed(16'sh0) : $signed(_GEN_328); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_624 = _T_69 ? $signed(16'sh0) : $signed(_GEN_329); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_625 = _T_69 ? $signed(16'sh0) : $signed(_GEN_330); // @[Conditional.scala 39:67 switch.scala 35:19]
  wire [15:0] _GEN_626 = _T_69 ? $signed(16'sh0) : $signed(_GEN_331); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_627 = _T_69 ? $signed(16'sh0) : $signed(_GEN_332); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_628 = _T_69 ? $signed(16'sh0) : $signed(_GEN_333); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_629 = _T_69 ? $signed(16'sh0) : $signed(_GEN_334); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_630 = _T_69 ? $signed(16'sh0) : $signed(_GEN_335); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_631 = _T_69 ? $signed(16'sh0) : $signed(_GEN_336); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_632 = _T_69 ? $signed(16'sh0) : $signed(_GEN_337); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_633 = _T_69 ? $signed(16'sh0) : $signed(_GEN_338); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_634 = _T_69 ? $signed(16'sh0) : $signed(_GEN_339); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_635 = _T_69 ? $signed(16'sh0) : $signed(_GEN_340); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_636 = _T_69 ? $signed(16'sh0) : $signed(_GEN_341); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_637 = _T_69 ? $signed(16'sh0) : $signed(_GEN_342); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_638 = _T_69 ? $signed(16'sh0) : $signed(_GEN_343); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_639 = _T_69 ? $signed(16'sh0) : $signed(_GEN_344); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_640 = _T_69 ? $signed(16'sh0) : $signed(_GEN_345); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_641 = _T_69 ? $signed(16'sh0) : $signed(_GEN_346); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_642 = _T_69 ? $signed(16'sh0) : $signed(_GEN_347); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_643 = _T_69 ? $signed(16'sh0) : $signed(_GEN_348); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_644 = _T_69 ? $signed(16'sh0) : $signed(_GEN_349); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_645 = _T_69 ? $signed(16'sh0) : $signed(_GEN_350); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_646 = _T_69 ? $signed(16'sh0) : $signed(_GEN_351); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_647 = _T_69 ? $signed(16'sh0) : $signed(_GEN_352); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_648 = _T_69 ? $signed(16'sh0) : $signed(_GEN_353); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_649 = _T_69 ? $signed(16'sh0) : $signed(_GEN_354); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_650 = _T_69 ? $signed(16'sh0) : $signed(_GEN_355); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_651 = _T_69 ? $signed(16'sh0) : $signed(_GEN_356); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_652 = _T_69 ? $signed(16'sh0) : $signed(_GEN_357); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_653 = _T_69 ? $signed(16'sh0) : $signed(_GEN_358); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_654 = _T_69 ? $signed(16'sh0) : $signed(_GEN_359); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_655 = _T_69 ? $signed(16'sh0) : $signed(_GEN_360); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_656 = _T_69 ? $signed(16'sh0) : $signed(_GEN_361); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_657 = _T_69 ? $signed(16'sh0) : $signed(_GEN_362); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_658 = _T_69 ? $signed(16'sh0) : $signed(_GEN_363); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_659 = _T_69 ? $signed(16'sh0) : $signed(_GEN_364); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_660 = _T_69 ? $signed(16'sh0) : $signed(_GEN_365); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_661 = _T_69 ? $signed(16'sh0) : $signed(_GEN_366); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_662 = _T_69 ? $signed(16'sh0) : $signed(_GEN_367); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_663 = _T_69 ? $signed(16'sh0) : $signed(_GEN_368); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_664 = _T_69 ? $signed(16'sh0) : $signed(_GEN_369); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_665 = _T_69 ? $signed(16'sh0) : $signed(_GEN_370); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_666 = _T_69 ? $signed(16'sh0) : $signed(_GEN_371); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_667 = _T_69 ? $signed(16'sh0) : $signed(_GEN_372); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_668 = _T_69 ? $signed(16'sh0) : $signed(_GEN_373); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_669 = _T_69 ? $signed(16'sh0) : $signed(_GEN_374); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_670 = _T_69 ? $signed(16'sh0) : $signed(_GEN_375); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_671 = _T_69 ? $signed(16'sh0) : $signed(_GEN_376); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_672 = _T_69 ? $signed(16'sh0) : $signed(_GEN_377); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_673 = _T_69 ? $signed(16'sh0) : $signed(_GEN_378); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_674 = _T_69 ? $signed(16'sh0) : $signed(_GEN_379); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_675 = _T_69 ? $signed(16'sh0) : $signed(_GEN_380); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_676 = _T_69 ? $signed(16'sh0) : $signed(_GEN_381); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_677 = _T_69 ? $signed(16'sh0) : $signed(_GEN_382); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_678 = _T_69 ? $signed(16'sh0) : $signed(_GEN_383); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_679 = _T_69 ? $signed(16'sh0) : $signed(_GEN_384); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_680 = _T_69 ? $signed(16'sh0) : $signed(_GEN_385); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_681 = _T_69 ? $signed(16'sh0) : $signed(_GEN_386); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_682 = _T_69 ? $signed(16'sh0) : $signed(_GEN_387); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_683 = _T_69 ? $signed(16'sh0) : $signed(_GEN_388); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_684 = _T_69 ? $signed(16'sh0) : $signed(_GEN_389); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_685 = _T_69 ? $signed(16'sh0) : $signed(_GEN_390); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_686 = _T_69 ? $signed(16'sh0) : $signed(_GEN_391); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_687 = _T_69 ? $signed(16'sh0) : $signed(_GEN_392); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_688 = _T_69 ? $signed(16'sh0) : $signed(_GEN_393); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_689 = _T_69 ? $signed(16'sh0) : $signed(_GEN_394); // @[Conditional.scala 39:67 switch.scala 36:18]
  wire [15:0] _GEN_690 = _T_69 ? $signed(cache_0) : $signed(_GEN_395); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_691 = _T_69 ? $signed(cache_1) : $signed(_GEN_396); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_692 = _T_69 ? $signed(cache_2) : $signed(_GEN_397); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_693 = _T_69 ? $signed(cache_3) : $signed(_GEN_398); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_694 = _T_69 ? $signed(cache_4) : $signed(_GEN_399); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_695 = _T_69 ? $signed(cache_5) : $signed(_GEN_400); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_696 = _T_69 ? $signed(cache_6) : $signed(_GEN_401); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_697 = _T_69 ? $signed(cache_7) : $signed(_GEN_402); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_698 = _T_69 ? $signed(cache_8) : $signed(_GEN_403); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_699 = _T_69 ? $signed(cache_9) : $signed(_GEN_404); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_700 = _T_69 ? $signed(cache_10) : $signed(_GEN_405); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_701 = _T_69 ? $signed(cache_11) : $signed(_GEN_406); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_702 = _T_69 ? $signed(cache_12) : $signed(_GEN_407); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_703 = _T_69 ? $signed(cache_13) : $signed(_GEN_408); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_704 = _T_69 ? $signed(cache_14) : $signed(_GEN_409); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_705 = _T_69 ? $signed(cache_15) : $signed(_GEN_410); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_706 = _T_69 ? $signed(cache_16) : $signed(_GEN_411); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_707 = _T_69 ? $signed(cache_17) : $signed(_GEN_412); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_708 = _T_69 ? $signed(cache_18) : $signed(_GEN_413); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_709 = _T_69 ? $signed(cache_19) : $signed(_GEN_414); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_710 = _T_69 ? $signed(cache_20) : $signed(_GEN_415); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_711 = _T_69 ? $signed(cache_21) : $signed(_GEN_416); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_712 = _T_69 ? $signed(cache_22) : $signed(_GEN_417); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_713 = _T_69 ? $signed(cache_23) : $signed(_GEN_418); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_714 = _T_69 ? $signed(cache_24) : $signed(_GEN_419); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_715 = _T_69 ? $signed(cache_25) : $signed(_GEN_420); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_716 = _T_69 ? $signed(cache_26) : $signed(_GEN_421); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_717 = _T_69 ? $signed(cache_27) : $signed(_GEN_422); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_718 = _T_69 ? $signed(cache_28) : $signed(_GEN_423); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_719 = _T_69 ? $signed(cache_29) : $signed(_GEN_424); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_720 = _T_69 ? $signed(cache_30) : $signed(_GEN_425); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_721 = _T_69 ? $signed(cache_31) : $signed(_GEN_426); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_722 = _T_69 ? $signed(cache_32) : $signed(_GEN_427); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_723 = _T_69 ? $signed(cache_33) : $signed(_GEN_428); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_724 = _T_69 ? $signed(cache_34) : $signed(_GEN_429); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_725 = _T_69 ? $signed(cache_35) : $signed(_GEN_430); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_726 = _T_69 ? $signed(cache_36) : $signed(_GEN_431); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_727 = _T_69 ? $signed(cache_37) : $signed(_GEN_432); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_728 = _T_69 ? $signed(cache_38) : $signed(_GEN_433); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_729 = _T_69 ? $signed(cache_39) : $signed(_GEN_434); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_730 = _T_69 ? $signed(cache_40) : $signed(_GEN_435); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_731 = _T_69 ? $signed(cache_41) : $signed(_GEN_436); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_732 = _T_69 ? $signed(cache_42) : $signed(_GEN_437); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_733 = _T_69 ? $signed(cache_43) : $signed(_GEN_438); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_734 = _T_69 ? $signed(cache_44) : $signed(_GEN_439); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_735 = _T_69 ? $signed(cache_45) : $signed(_GEN_440); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_736 = _T_69 ? $signed(cache_46) : $signed(_GEN_441); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_737 = _T_69 ? $signed(cache_47) : $signed(_GEN_442); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_738 = _T_69 ? $signed(cache_48) : $signed(_GEN_443); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_739 = _T_69 ? $signed(cache_49) : $signed(_GEN_444); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_740 = _T_69 ? $signed(cache_50) : $signed(_GEN_445); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_741 = _T_69 ? $signed(cache_51) : $signed(_GEN_446); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_742 = _T_69 ? $signed(cache_52) : $signed(_GEN_447); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_743 = _T_69 ? $signed(cache_53) : $signed(_GEN_448); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_744 = _T_69 ? $signed(cache_54) : $signed(_GEN_449); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_745 = _T_69 ? $signed(cache_55) : $signed(_GEN_450); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_746 = _T_69 ? $signed(cache_56) : $signed(_GEN_451); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_747 = _T_69 ? $signed(cache_57) : $signed(_GEN_452); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_748 = _T_69 ? $signed(cache_58) : $signed(_GEN_453); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_749 = _T_69 ? $signed(cache_59) : $signed(_GEN_454); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_750 = _T_69 ? $signed(cache_60) : $signed(_GEN_455); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_751 = _T_69 ? $signed(cache_61) : $signed(_GEN_456); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_752 = _T_69 ? $signed(cache_62) : $signed(_GEN_457); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_753 = _T_69 ? $signed(cache_63) : $signed(_GEN_458); // @[Conditional.scala 39:67 switch.scala 30:24]
  wire [15:0] _GEN_754 = _T_66 ? $signed(io_from_right_0) : $signed(_GEN_526); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_755 = _T_66 ? $signed(io_from_right_1) : $signed(_GEN_527); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_756 = _T_66 ? $signed(io_from_right_2) : $signed(_GEN_528); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_757 = _T_66 ? $signed(io_from_right_3) : $signed(_GEN_529); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_758 = _T_66 ? $signed(io_from_right_4) : $signed(_GEN_530); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_759 = _T_66 ? $signed(io_from_right_5) : $signed(_GEN_531); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_760 = _T_66 ? $signed(io_from_right_6) : $signed(_GEN_532); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_761 = _T_66 ? $signed(io_from_right_7) : $signed(_GEN_533); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_762 = _T_66 ? $signed(io_from_left_0) : $signed(_GEN_534); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_763 = _T_66 ? $signed(io_from_left_1) : $signed(_GEN_535); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_764 = _T_66 ? $signed(io_from_left_2) : $signed(_GEN_536); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_765 = _T_66 ? $signed(io_from_left_3) : $signed(_GEN_537); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_766 = _T_66 ? $signed(io_from_left_4) : $signed(_GEN_538); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_767 = _T_66 ? $signed(io_from_left_5) : $signed(_GEN_539); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_768 = _T_66 ? $signed(io_from_left_6) : $signed(_GEN_540); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_769 = _T_66 ? $signed(io_from_left_7) : $signed(_GEN_541); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_770 = _T_66 ? $signed(io_from_down_0) : $signed(_GEN_542); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_771 = _T_66 ? $signed(io_from_down_1) : $signed(_GEN_543); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_772 = _T_66 ? $signed(io_from_down_2) : $signed(_GEN_544); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_773 = _T_66 ? $signed(io_from_down_3) : $signed(_GEN_545); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_774 = _T_66 ? $signed(io_from_down_4) : $signed(_GEN_546); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_775 = _T_66 ? $signed(io_from_down_5) : $signed(_GEN_547); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_776 = _T_66 ? $signed(io_from_down_6) : $signed(_GEN_548); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_777 = _T_66 ? $signed(io_from_down_7) : $signed(_GEN_549); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_778 = _T_66 ? $signed(io_from_down_8) : $signed(_GEN_550); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_779 = _T_66 ? $signed(io_from_down_9) : $signed(_GEN_551); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_780 = _T_66 ? $signed(io_from_up_0) : $signed(_GEN_552); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_781 = _T_66 ? $signed(io_from_up_1) : $signed(_GEN_553); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_782 = _T_66 ? $signed(io_from_up_2) : $signed(_GEN_554); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_783 = _T_66 ? $signed(io_from_up_3) : $signed(_GEN_555); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_784 = _T_66 ? $signed(io_from_up_4) : $signed(_GEN_556); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_785 = _T_66 ? $signed(io_from_up_5) : $signed(_GEN_557); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_786 = _T_66 ? $signed(io_from_up_6) : $signed(_GEN_558); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_787 = _T_66 ? $signed(io_from_up_7) : $signed(_GEN_559); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_788 = _T_66 ? $signed(io_from_up_8) : $signed(_GEN_560); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_789 = _T_66 ? $signed(io_from_up_9) : $signed(_GEN_561); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_790 = _T_66 ? $signed(io_from_mat_0) : $signed(_GEN_562); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_791 = _T_66 ? $signed(io_from_mat_1) : $signed(_GEN_563); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_792 = _T_66 ? $signed(io_from_mat_2) : $signed(_GEN_564); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_793 = _T_66 ? $signed(io_from_mat_3) : $signed(_GEN_565); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_794 = _T_66 ? $signed(io_from_mat_4) : $signed(_GEN_566); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_795 = _T_66 ? $signed(io_from_mat_5) : $signed(_GEN_567); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_796 = _T_66 ? $signed(io_from_mat_6) : $signed(_GEN_568); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_797 = _T_66 ? $signed(io_from_mat_7) : $signed(_GEN_569); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_798 = _T_66 ? $signed(io_from_mat_8) : $signed(_GEN_570); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_799 = _T_66 ? $signed(io_from_mat_9) : $signed(_GEN_571); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_800 = _T_66 ? $signed(io_from_mat_10) : $signed(_GEN_572); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_801 = _T_66 ? $signed(io_from_mat_11) : $signed(_GEN_573); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_802 = _T_66 ? $signed(io_from_mat_12) : $signed(_GEN_574); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_803 = _T_66 ? $signed(io_from_mat_13) : $signed(_GEN_575); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_804 = _T_66 ? $signed(io_from_mat_14) : $signed(_GEN_576); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_805 = _T_66 ? $signed(io_from_mat_15) : $signed(_GEN_577); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_806 = _T_66 ? $signed(io_from_mat_16) : $signed(_GEN_578); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_807 = _T_66 ? $signed(io_from_mat_17) : $signed(_GEN_579); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_808 = _T_66 ? $signed(io_from_mat_18) : $signed(_GEN_580); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_809 = _T_66 ? $signed(io_from_mat_19) : $signed(_GEN_581); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_810 = _T_66 ? $signed(io_from_mat_20) : $signed(_GEN_582); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_811 = _T_66 ? $signed(io_from_mat_21) : $signed(_GEN_583); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_812 = _T_66 ? $signed(io_from_mat_22) : $signed(_GEN_584); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_813 = _T_66 ? $signed(io_from_mat_23) : $signed(_GEN_585); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_814 = _T_66 ? $signed(io_from_mat_24) : $signed(_GEN_586); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_815 = _T_66 ? $signed(io_from_mat_25) : $signed(_GEN_587); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_816 = _T_66 ? $signed(io_from_mat_26) : $signed(_GEN_588); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_817 = _T_66 ? $signed(io_from_mat_27) : $signed(_GEN_589); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_818 = _T_66 ? $signed(io_from_mat_28) : $signed(_GEN_590); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_819 = _T_66 ? $signed(io_from_mat_29) : $signed(_GEN_591); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_820 = _T_66 ? $signed(io_from_mat_30) : $signed(_GEN_592); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_821 = _T_66 ? $signed(io_from_mat_31) : $signed(_GEN_593); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_822 = _T_66 ? $signed(io_from_mat_32) : $signed(_GEN_594); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_823 = _T_66 ? $signed(io_from_mat_33) : $signed(_GEN_595); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_824 = _T_66 ? $signed(io_from_mat_34) : $signed(_GEN_596); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_825 = _T_66 ? $signed(io_from_mat_35) : $signed(_GEN_597); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_826 = _T_66 ? $signed(io_from_mat_36) : $signed(_GEN_598); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_827 = _T_66 ? $signed(io_from_mat_37) : $signed(_GEN_599); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_828 = _T_66 ? $signed(io_from_mat_38) : $signed(_GEN_600); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_829 = _T_66 ? $signed(io_from_mat_39) : $signed(_GEN_601); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_830 = _T_66 ? $signed(io_from_mat_40) : $signed(_GEN_602); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_831 = _T_66 ? $signed(io_from_mat_41) : $signed(_GEN_603); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_832 = _T_66 ? $signed(io_from_mat_42) : $signed(_GEN_604); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_833 = _T_66 ? $signed(io_from_mat_43) : $signed(_GEN_605); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_834 = _T_66 ? $signed(io_from_mat_44) : $signed(_GEN_606); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_835 = _T_66 ? $signed(io_from_mat_45) : $signed(_GEN_607); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_836 = _T_66 ? $signed(io_from_mat_46) : $signed(_GEN_608); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_837 = _T_66 ? $signed(io_from_mat_47) : $signed(_GEN_609); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_838 = _T_66 ? $signed(io_from_mat_48) : $signed(_GEN_610); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_839 = _T_66 ? $signed(io_from_mat_49) : $signed(_GEN_611); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_840 = _T_66 ? $signed(io_from_mat_50) : $signed(_GEN_612); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_841 = _T_66 ? $signed(io_from_mat_51) : $signed(_GEN_613); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_842 = _T_66 ? $signed(io_from_mat_52) : $signed(_GEN_614); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_843 = _T_66 ? $signed(io_from_mat_53) : $signed(_GEN_615); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_844 = _T_66 ? $signed(io_from_mat_54) : $signed(_GEN_616); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_845 = _T_66 ? $signed(io_from_mat_55) : $signed(_GEN_617); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_846 = _T_66 ? $signed(io_from_mat_56) : $signed(_GEN_618); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_847 = _T_66 ? $signed(io_from_mat_57) : $signed(_GEN_619); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_848 = _T_66 ? $signed(io_from_mat_58) : $signed(_GEN_620); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_849 = _T_66 ? $signed(io_from_mat_59) : $signed(_GEN_621); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_850 = _T_66 ? $signed(io_from_mat_60) : $signed(_GEN_622); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_851 = _T_66 ? $signed(io_from_mat_61) : $signed(_GEN_623); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_852 = _T_66 ? $signed(io_from_mat_62) : $signed(_GEN_624); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_853 = _T_66 ? $signed(io_from_mat_63) : $signed(_GEN_625); // @[Conditional.scala 40:58 switch.scala 45:31]
  wire [15:0] _GEN_854 = _T_66 ? $signed(io_from_weight_0) : $signed(_GEN_626); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire [15:0] _GEN_855 = _T_66 ? $signed(io_from_weight_1) : $signed(_GEN_627); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire [15:0] _GEN_856 = _T_66 ? $signed(io_from_weight_2) : $signed(_GEN_628); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire [15:0] _GEN_857 = _T_66 ? $signed(io_from_weight_3) : $signed(_GEN_629); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire [15:0] _GEN_858 = _T_66 ? $signed(io_from_weight_4) : $signed(_GEN_630); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire [15:0] _GEN_859 = _T_66 ? $signed(io_from_weight_5) : $signed(_GEN_631); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire [15:0] _GEN_860 = _T_66 ? $signed(io_from_weight_6) : $signed(_GEN_632); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire [15:0] _GEN_861 = _T_66 ? $signed(io_from_weight_7) : $signed(_GEN_633); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire [15:0] _GEN_862 = _T_66 ? $signed(io_from_weight_8) : $signed(_GEN_634); // @[Conditional.scala 40:58 switch.scala 47:45]
  wire  _GEN_863 = _T_66 | _GEN_525; // @[Conditional.scala 40:58 switch.scala 48:38]
  wire [15:0] _GEN_930 = _T_66 ? $signed(16'sh0) : $signed(_GEN_635); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_931 = _T_66 ? $signed(16'sh0) : $signed(_GEN_636); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_932 = _T_66 ? $signed(16'sh0) : $signed(_GEN_637); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_933 = _T_66 ? $signed(16'sh0) : $signed(_GEN_638); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_934 = _T_66 ? $signed(16'sh0) : $signed(_GEN_639); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_935 = _T_66 ? $signed(16'sh0) : $signed(_GEN_640); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_936 = _T_66 ? $signed(16'sh0) : $signed(_GEN_641); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_937 = _T_66 ? $signed(16'sh0) : $signed(_GEN_642); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_938 = _T_66 ? $signed(16'sh0) : $signed(_GEN_643); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_939 = _T_66 ? $signed(16'sh0) : $signed(_GEN_644); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_940 = _T_66 ? $signed(16'sh0) : $signed(_GEN_645); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_941 = _T_66 ? $signed(16'sh0) : $signed(_GEN_646); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_942 = _T_66 ? $signed(16'sh0) : $signed(_GEN_647); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_943 = _T_66 ? $signed(16'sh0) : $signed(_GEN_648); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_944 = _T_66 ? $signed(16'sh0) : $signed(_GEN_649); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_945 = _T_66 ? $signed(16'sh0) : $signed(_GEN_650); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_946 = _T_66 ? $signed(16'sh0) : $signed(_GEN_651); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_947 = _T_66 ? $signed(16'sh0) : $signed(_GEN_652); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_948 = _T_66 ? $signed(16'sh0) : $signed(_GEN_653); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_949 = _T_66 ? $signed(16'sh0) : $signed(_GEN_654); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_950 = _T_66 ? $signed(16'sh0) : $signed(_GEN_655); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_951 = _T_66 ? $signed(16'sh0) : $signed(_GEN_656); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_952 = _T_66 ? $signed(16'sh0) : $signed(_GEN_657); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_953 = _T_66 ? $signed(16'sh0) : $signed(_GEN_658); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_954 = _T_66 ? $signed(16'sh0) : $signed(_GEN_659); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_955 = _T_66 ? $signed(16'sh0) : $signed(_GEN_660); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_956 = _T_66 ? $signed(16'sh0) : $signed(_GEN_661); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_957 = _T_66 ? $signed(16'sh0) : $signed(_GEN_662); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_958 = _T_66 ? $signed(16'sh0) : $signed(_GEN_663); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_959 = _T_66 ? $signed(16'sh0) : $signed(_GEN_664); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_960 = _T_66 ? $signed(16'sh0) : $signed(_GEN_665); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_961 = _T_66 ? $signed(16'sh0) : $signed(_GEN_666); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_962 = _T_66 ? $signed(16'sh0) : $signed(_GEN_667); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_963 = _T_66 ? $signed(16'sh0) : $signed(_GEN_668); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_964 = _T_66 ? $signed(16'sh0) : $signed(_GEN_669); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_965 = _T_66 ? $signed(16'sh0) : $signed(_GEN_670); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_966 = _T_66 ? $signed(16'sh0) : $signed(_GEN_671); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_967 = _T_66 ? $signed(16'sh0) : $signed(_GEN_672); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_968 = _T_66 ? $signed(16'sh0) : $signed(_GEN_673); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_969 = _T_66 ? $signed(16'sh0) : $signed(_GEN_674); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_970 = _T_66 ? $signed(16'sh0) : $signed(_GEN_675); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_971 = _T_66 ? $signed(16'sh0) : $signed(_GEN_676); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_972 = _T_66 ? $signed(16'sh0) : $signed(_GEN_677); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_973 = _T_66 ? $signed(16'sh0) : $signed(_GEN_678); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_974 = _T_66 ? $signed(16'sh0) : $signed(_GEN_679); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_975 = _T_66 ? $signed(16'sh0) : $signed(_GEN_680); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_976 = _T_66 ? $signed(16'sh0) : $signed(_GEN_681); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_977 = _T_66 ? $signed(16'sh0) : $signed(_GEN_682); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_978 = _T_66 ? $signed(16'sh0) : $signed(_GEN_683); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_979 = _T_66 ? $signed(16'sh0) : $signed(_GEN_684); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_980 = _T_66 ? $signed(16'sh0) : $signed(_GEN_685); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_981 = _T_66 ? $signed(16'sh0) : $signed(_GEN_686); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_982 = _T_66 ? $signed(16'sh0) : $signed(_GEN_687); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_983 = _T_66 ? $signed(16'sh0) : $signed(_GEN_688); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_984 = _T_66 ? $signed(16'sh0) : $signed(_GEN_689); // @[Conditional.scala 40:58 switch.scala 36:18]
  wire [15:0] _GEN_1049 = io_valid_in ? $signed(_GEN_754) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1050 = io_valid_in ? $signed(_GEN_755) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1051 = io_valid_in ? $signed(_GEN_756) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1052 = io_valid_in ? $signed(_GEN_757) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1053 = io_valid_in ? $signed(_GEN_758) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1054 = io_valid_in ? $signed(_GEN_759) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1055 = io_valid_in ? $signed(_GEN_760) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1056 = io_valid_in ? $signed(_GEN_761) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1057 = io_valid_in ? $signed(_GEN_762) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1058 = io_valid_in ? $signed(_GEN_763) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1059 = io_valid_in ? $signed(_GEN_764) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1060 = io_valid_in ? $signed(_GEN_765) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1061 = io_valid_in ? $signed(_GEN_766) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1062 = io_valid_in ? $signed(_GEN_767) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1063 = io_valid_in ? $signed(_GEN_768) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1064 = io_valid_in ? $signed(_GEN_769) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1065 = io_valid_in ? $signed(_GEN_770) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1066 = io_valid_in ? $signed(_GEN_771) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1067 = io_valid_in ? $signed(_GEN_772) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1068 = io_valid_in ? $signed(_GEN_773) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1069 = io_valid_in ? $signed(_GEN_774) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1070 = io_valid_in ? $signed(_GEN_775) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1071 = io_valid_in ? $signed(_GEN_776) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1072 = io_valid_in ? $signed(_GEN_777) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1073 = io_valid_in ? $signed(_GEN_778) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1074 = io_valid_in ? $signed(_GEN_779) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1075 = io_valid_in ? $signed(_GEN_780) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1076 = io_valid_in ? $signed(_GEN_781) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1077 = io_valid_in ? $signed(_GEN_782) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1078 = io_valid_in ? $signed(_GEN_783) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1079 = io_valid_in ? $signed(_GEN_784) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1080 = io_valid_in ? $signed(_GEN_785) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1081 = io_valid_in ? $signed(_GEN_786) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1082 = io_valid_in ? $signed(_GEN_787) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1083 = io_valid_in ? $signed(_GEN_788) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1084 = io_valid_in ? $signed(_GEN_789) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1085 = io_valid_in ? $signed(_GEN_790) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1086 = io_valid_in ? $signed(_GEN_791) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1087 = io_valid_in ? $signed(_GEN_792) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1088 = io_valid_in ? $signed(_GEN_793) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1089 = io_valid_in ? $signed(_GEN_794) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1090 = io_valid_in ? $signed(_GEN_795) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1091 = io_valid_in ? $signed(_GEN_796) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1092 = io_valid_in ? $signed(_GEN_797) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1093 = io_valid_in ? $signed(_GEN_798) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1094 = io_valid_in ? $signed(_GEN_799) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1095 = io_valid_in ? $signed(_GEN_800) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1096 = io_valid_in ? $signed(_GEN_801) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1097 = io_valid_in ? $signed(_GEN_802) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1098 = io_valid_in ? $signed(_GEN_803) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1099 = io_valid_in ? $signed(_GEN_804) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1100 = io_valid_in ? $signed(_GEN_805) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1101 = io_valid_in ? $signed(_GEN_806) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1102 = io_valid_in ? $signed(_GEN_807) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1103 = io_valid_in ? $signed(_GEN_808) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1104 = io_valid_in ? $signed(_GEN_809) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1105 = io_valid_in ? $signed(_GEN_810) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1106 = io_valid_in ? $signed(_GEN_811) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1107 = io_valid_in ? $signed(_GEN_812) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1108 = io_valid_in ? $signed(_GEN_813) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1109 = io_valid_in ? $signed(_GEN_814) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1110 = io_valid_in ? $signed(_GEN_815) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1111 = io_valid_in ? $signed(_GEN_816) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1112 = io_valid_in ? $signed(_GEN_817) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1113 = io_valid_in ? $signed(_GEN_818) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1114 = io_valid_in ? $signed(_GEN_819) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1115 = io_valid_in ? $signed(_GEN_820) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1116 = io_valid_in ? $signed(_GEN_821) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1117 = io_valid_in ? $signed(_GEN_822) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1118 = io_valid_in ? $signed(_GEN_823) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1119 = io_valid_in ? $signed(_GEN_824) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1120 = io_valid_in ? $signed(_GEN_825) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1121 = io_valid_in ? $signed(_GEN_826) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1122 = io_valid_in ? $signed(_GEN_827) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1123 = io_valid_in ? $signed(_GEN_828) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1124 = io_valid_in ? $signed(_GEN_829) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1125 = io_valid_in ? $signed(_GEN_830) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1126 = io_valid_in ? $signed(_GEN_831) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1127 = io_valid_in ? $signed(_GEN_832) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1128 = io_valid_in ? $signed(_GEN_833) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1129 = io_valid_in ? $signed(_GEN_834) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1130 = io_valid_in ? $signed(_GEN_835) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1131 = io_valid_in ? $signed(_GEN_836) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1132 = io_valid_in ? $signed(_GEN_837) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1133 = io_valid_in ? $signed(_GEN_838) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1134 = io_valid_in ? $signed(_GEN_839) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1135 = io_valid_in ? $signed(_GEN_840) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1136 = io_valid_in ? $signed(_GEN_841) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1137 = io_valid_in ? $signed(_GEN_842) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1138 = io_valid_in ? $signed(_GEN_843) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1139 = io_valid_in ? $signed(_GEN_844) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1140 = io_valid_in ? $signed(_GEN_845) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1141 = io_valid_in ? $signed(_GEN_846) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1142 = io_valid_in ? $signed(_GEN_847) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1143 = io_valid_in ? $signed(_GEN_848) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1144 = io_valid_in ? $signed(_GEN_849) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1145 = io_valid_in ? $signed(_GEN_850) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1146 = io_valid_in ? $signed(_GEN_851) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1147 = io_valid_in ? $signed(_GEN_852) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1148 = io_valid_in ? $signed(_GEN_853) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 35:19]
  wire [15:0] _GEN_1149 = io_valid_in ? $signed(_GEN_854) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1150 = io_valid_in ? $signed(_GEN_855) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1151 = io_valid_in ? $signed(_GEN_856) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1152 = io_valid_in ? $signed(_GEN_857) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1153 = io_valid_in ? $signed(_GEN_858) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1154 = io_valid_in ? $signed(_GEN_859) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1155 = io_valid_in ? $signed(_GEN_860) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1156 = io_valid_in ? $signed(_GEN_861) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1157 = io_valid_in ? $signed(_GEN_862) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire  _GEN_1158 = io_valid_in & _GEN_863; // @[switch.scala 42:28 switch.scala 33:26]
  wire [15:0] _GEN_1225 = io_valid_in ? $signed(_GEN_930) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1226 = io_valid_in ? $signed(_GEN_931) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1227 = io_valid_in ? $signed(_GEN_932) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1228 = io_valid_in ? $signed(_GEN_933) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1229 = io_valid_in ? $signed(_GEN_934) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1230 = io_valid_in ? $signed(_GEN_935) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1231 = io_valid_in ? $signed(_GEN_936) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1232 = io_valid_in ? $signed(_GEN_937) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1233 = io_valid_in ? $signed(_GEN_938) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1234 = io_valid_in ? $signed(_GEN_939) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1235 = io_valid_in ? $signed(_GEN_940) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1236 = io_valid_in ? $signed(_GEN_941) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1237 = io_valid_in ? $signed(_GEN_942) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1238 = io_valid_in ? $signed(_GEN_943) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1239 = io_valid_in ? $signed(_GEN_944) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1240 = io_valid_in ? $signed(_GEN_945) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1241 = io_valid_in ? $signed(_GEN_946) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1242 = io_valid_in ? $signed(_GEN_947) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1243 = io_valid_in ? $signed(_GEN_948) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1244 = io_valid_in ? $signed(_GEN_949) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1245 = io_valid_in ? $signed(_GEN_950) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1246 = io_valid_in ? $signed(_GEN_951) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1247 = io_valid_in ? $signed(_GEN_952) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1248 = io_valid_in ? $signed(_GEN_953) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1249 = io_valid_in ? $signed(_GEN_954) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1250 = io_valid_in ? $signed(_GEN_955) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1251 = io_valid_in ? $signed(_GEN_956) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1252 = io_valid_in ? $signed(_GEN_957) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1253 = io_valid_in ? $signed(_GEN_958) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1254 = io_valid_in ? $signed(_GEN_959) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1255 = io_valid_in ? $signed(_GEN_960) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1256 = io_valid_in ? $signed(_GEN_961) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1257 = io_valid_in ? $signed(_GEN_962) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1258 = io_valid_in ? $signed(_GEN_963) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1259 = io_valid_in ? $signed(_GEN_964) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1260 = io_valid_in ? $signed(_GEN_965) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1261 = io_valid_in ? $signed(_GEN_966) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1262 = io_valid_in ? $signed(_GEN_967) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1263 = io_valid_in ? $signed(_GEN_968) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1264 = io_valid_in ? $signed(_GEN_969) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1265 = io_valid_in ? $signed(_GEN_970) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1266 = io_valid_in ? $signed(_GEN_971) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1267 = io_valid_in ? $signed(_GEN_972) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1268 = io_valid_in ? $signed(_GEN_973) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1269 = io_valid_in ? $signed(_GEN_974) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1270 = io_valid_in ? $signed(_GEN_975) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1271 = io_valid_in ? $signed(_GEN_976) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1272 = io_valid_in ? $signed(_GEN_977) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1273 = io_valid_in ? $signed(_GEN_978) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1274 = io_valid_in ? $signed(_GEN_979) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1275 = io_valid_in ? $signed(_GEN_980) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1276 = io_valid_in ? $signed(_GEN_981) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1277 = io_valid_in ? $signed(_GEN_982) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1278 = io_valid_in ? $signed(_GEN_983) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire [15:0] _GEN_1279 = io_valid_in ? $signed(_GEN_984) : $signed(16'sh0); // @[switch.scala 42:28 switch.scala 36:18]
  wire  _GEN_1345 = io_flag_job | state_cend; // @[switch.scala 39:22 utils.scala 22:14 switch.scala 31:24]
  assign io_valid_out_calc8x8 = io_flag_job ? 1'h0 : _GEN_1158; // @[switch.scala 39:22 switch.scala 33:26]
  assign io_to_calc8x8_mat_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1085); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1086); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1087); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1088); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1089); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1090); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1091); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1092); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1093); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1094); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_10 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1095); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_11 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1096); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_12 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1097); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_13 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1098); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_14 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1099); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_15 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1100); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_16 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1101); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_17 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1102); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_18 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1103); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_19 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1104); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_20 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1105); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_21 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1106); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_22 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1107); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_23 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1108); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_24 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1109); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_25 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1110); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_26 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1111); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_27 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1112); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_28 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1113); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_29 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1114); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_30 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1115); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_31 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1116); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_32 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1117); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_33 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1118); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_34 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1119); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_35 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1120); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_36 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1121); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_37 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1122); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_38 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1123); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_39 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1124); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_40 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1125); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_41 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1126); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_42 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1127); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_43 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1128); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_44 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1129); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_45 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1130); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_46 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1131); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_47 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1132); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_48 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1133); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_49 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1134); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_50 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1135); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_51 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1136); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_52 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1137); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_53 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1138); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_54 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1139); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_55 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1140); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_56 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1141); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_57 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1142); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_58 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1143); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_59 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1144); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_60 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1145); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_61 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1146); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_62 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1147); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_mat_63 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1148); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1075); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1076); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1077); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1078); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1079); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1080); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1081); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1082); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1083); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_up_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1084); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1065); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1066); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1067); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1068); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1069); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1070); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1071); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1072); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1073); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_down_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1074); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_left_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1057); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_left_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1058); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_left_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1059); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_left_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1060); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_left_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1061); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_left_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1062); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_left_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1063); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_left_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1064); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_right_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1049); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_right_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1050); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_right_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1051); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_right_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1052); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_right_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1053); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_right_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1054); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_right_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1055); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_calc8x8_right_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1056); // @[switch.scala 39:22 switch.scala 35:19]
  assign io_to_weight_0_real_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1149); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1150); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1151); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1152); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1153); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1154); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1155); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1156); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1157); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1225); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_10 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1226); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_11 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1227); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_12 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1228); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_13 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1229); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_14 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1230); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_0_real_15 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1231); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1232); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1233); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1234); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1235); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1236); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1237); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1238); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1239); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1240); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1241); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_10 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1242); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_11 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1243); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_12 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1244); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_13 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1245); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_14 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1246); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_1_real_15 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1247); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1248); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1249); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1250); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1251); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1252); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1253); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1254); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1255); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1256); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1257); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_10 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1258); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_11 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1259); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_12 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1260); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_13 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1261); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_14 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1262); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_2_real_15 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1263); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_0 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1264); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_1 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1265); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_2 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1266); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_3 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1267); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_4 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1268); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_5 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1269); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_6 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1270); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_7 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1271); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_8 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1272); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_9 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1273); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_10 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1274); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_11 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1275); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_12 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1276); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_13 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1277); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_14 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1278); // @[switch.scala 39:22 switch.scala 36:18]
  assign io_to_weight_3_real_15 = io_flag_job ? $signed(16'sh0) : $signed(_GEN_1279); // @[switch.scala 39:22 switch.scala 36:18]
  always @(posedge clock) begin
    if (reset) begin // @[switch.scala 28:27]
      job_type <= 2'h0; // @[switch.scala 28:27]
    end else if (io_flag_job) begin // @[switch.scala 39:22]
      job_type <= io_job; // @[switch.scala 40:18]
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_0 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_0 <= _GEN_690;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_1 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_1 <= _GEN_691;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_2 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_2 <= _GEN_692;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_3 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_3 <= _GEN_693;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_4 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_4 <= _GEN_694;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_5 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_5 <= _GEN_695;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_6 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_6 <= _GEN_696;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_7 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_7 <= _GEN_697;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_8 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_8 <= _GEN_698;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_9 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_9 <= _GEN_699;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_10 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_10 <= _GEN_700;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_11 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_11 <= _GEN_701;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_12 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_12 <= _GEN_702;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_13 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_13 <= _GEN_703;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_14 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_14 <= _GEN_704;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_15 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_15 <= _GEN_705;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_16 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_16 <= _GEN_706;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_17 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_17 <= _GEN_707;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_18 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_18 <= _GEN_708;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_19 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_19 <= _GEN_709;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_20 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_20 <= _GEN_710;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_21 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_21 <= _GEN_711;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_22 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_22 <= _GEN_712;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_23 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_23 <= _GEN_713;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_24 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_24 <= _GEN_714;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_25 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_25 <= _GEN_715;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_26 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_26 <= _GEN_716;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_27 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_27 <= _GEN_717;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_28 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_28 <= _GEN_718;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_29 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_29 <= _GEN_719;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_30 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_30 <= _GEN_720;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_31 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_31 <= _GEN_721;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_32 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_32 <= _GEN_722;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_33 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_33 <= _GEN_723;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_34 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_34 <= _GEN_724;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_35 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_35 <= _GEN_725;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_36 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_36 <= _GEN_726;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_37 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_37 <= _GEN_727;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_38 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_38 <= _GEN_728;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_39 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_39 <= _GEN_729;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_40 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_40 <= _GEN_730;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_41 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_41 <= _GEN_731;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_42 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_42 <= _GEN_732;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_43 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_43 <= _GEN_733;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_44 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_44 <= _GEN_734;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_45 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_45 <= _GEN_735;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_46 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_46 <= _GEN_736;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_47 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_47 <= _GEN_737;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_48 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_48 <= _GEN_738;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_49 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_49 <= _GEN_739;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_50 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_50 <= _GEN_740;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_51 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_51 <= _GEN_741;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_52 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_52 <= _GEN_742;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_53 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_53 <= _GEN_743;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_54 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_54 <= _GEN_744;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_55 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_55 <= _GEN_745;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_56 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_56 <= _GEN_746;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_57 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_57 <= _GEN_747;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_58 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_58 <= _GEN_748;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_59 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_59 <= _GEN_749;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_60 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_60 <= _GEN_750;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_61 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_61 <= _GEN_751;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_62 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_62 <= _GEN_752;
        end
      end
    end
    if (reset) begin // @[switch.scala 30:24]
      cache_63 <= 16'sh0; // @[switch.scala 30:24]
    end else if (!(io_flag_job)) begin // @[switch.scala 39:22]
      if (io_valid_in) begin // @[switch.scala 42:28]
        if (!(_T_66)) begin // @[Conditional.scala 40:58]
          cache_63 <= _GEN_753;
        end
      end
    end
    if (reset) begin // @[switch.scala 31:24]
      state_ccnt <= 1'h0; // @[switch.scala 31:24]
    end else if (io_flag_job) begin // @[switch.scala 39:22]
      state_ccnt <= 1'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[switch.scala 42:28]
      if (!(_T_66)) begin // @[Conditional.scala 40:58]
        state_ccnt <= _GEN_524;
      end
    end
    if (reset) begin // @[switch.scala 31:24]
      state_cend <= 1'h0; // @[switch.scala 31:24]
    end else begin
      state_cend <= _GEN_1345;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  job_type = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cache_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  cache_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  cache_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  cache_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  cache_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  cache_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  cache_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  cache_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  cache_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  cache_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  cache_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  cache_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  cache_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  cache_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  cache_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  cache_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  cache_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  cache_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  cache_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  cache_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  cache_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  cache_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  cache_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  cache_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  cache_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  cache_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  cache_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  cache_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  cache_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  cache_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  cache_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  cache_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  cache_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  cache_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  cache_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  cache_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  cache_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  cache_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  cache_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  cache_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  cache_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  cache_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  cache_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  cache_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  cache_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  cache_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  cache_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  cache_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  cache_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  cache_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  cache_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  cache_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  cache_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  cache_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  cache_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  cache_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  cache_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  cache_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  cache_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  cache_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  cache_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  cache_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  cache_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  cache_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  state_ccnt = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  state_cend = _RAND_66[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WeightReader(
  input         clock,
  input         reset,
  input         io_valid_in,
  input         io_flag_job,
  input  [13:0] io_addr_end,
  output [13:0] io_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [13:0] now_addr_ccnt; // @[read_weight.scala 15:27]
  reg [13:0] now_addr_cend; // @[read_weight.scala 15:27]
  wire  nxt = now_addr_ccnt == now_addr_cend; // @[utils.scala 17:20]
  wire [13:0] _now_addr_ccnt_T_1 = now_addr_ccnt + 14'h1; // @[utils.scala 18:35]
  assign io_addr = now_addr_ccnt; // @[read_weight.scala 16:13]
  always @(posedge clock) begin
    if (reset) begin // @[read_weight.scala 15:27]
      now_addr_ccnt <= 14'h0; // @[read_weight.scala 15:27]
    end else if (io_flag_job) begin // @[read_weight.scala 18:22]
      now_addr_ccnt <= 14'h0; // @[utils.scala 27:14]
    end else if (io_valid_in) begin // @[read_weight.scala 20:28]
      if (nxt) begin // @[utils.scala 18:20]
        now_addr_ccnt <= 14'h0;
      end else begin
        now_addr_ccnt <= _now_addr_ccnt_T_1;
      end
    end
    if (reset) begin // @[read_weight.scala 15:27]
      now_addr_cend <= 14'h0; // @[read_weight.scala 15:27]
    end else if (io_flag_job) begin // @[read_weight.scala 18:22]
      now_addr_cend <= io_addr_end; // @[utils.scala 26:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  now_addr_ccnt = _RAND_0[13:0];
  _RAND_1 = {1{`RANDOM}};
  now_addr_cend = _RAND_1[13:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DSP48(
  input  [17:0] io_in_a,
  input  [24:0] io_in_b,
  output [42:0] io_out
);
  assign io_out = $signed(io_in_a) * $signed(io_in_b); // @[core.scala 53:22]
endmodule
module Core(
  input  [17:0] io_w_a,
  input  [24:0] io_in_b,
  input         io_flag,
  output [42:0] io_result
);
  wire [17:0] dsp48_io_in_a; // @[core.scala 21:23]
  wire [24:0] dsp48_io_in_b; // @[core.scala 21:23]
  wire [42:0] dsp48_io_out; // @[core.scala 21:23]
  wire  _T_2 = ~io_flag; // @[Conditional.scala 37:30]
  wire [15:0] _GEN_0 = io_in_b[24] ? $signed(16'sh7fff) : $signed(16'sh199a); // @[core.scala 27:30 core.scala 28:31 core.scala 30:31]
  wire [17:0] _GEN_1 = io_flag ? $signed(io_w_a) : $signed(18'sh0); // @[Conditional.scala 39:67 core.scala 34:27 core.scala 23:19]
  DSP48 dsp48 ( // @[core.scala 21:23]
    .io_in_a(dsp48_io_in_a),
    .io_in_b(dsp48_io_in_b),
    .io_out(dsp48_io_out)
  );
  assign io_result = dsp48_io_out; // @[core.scala 24:15]
  assign dsp48_io_in_a = _T_2 ? $signed({{2{_GEN_0[15]}},_GEN_0}) : $signed(_GEN_1); // @[Conditional.scala 40:58]
  assign dsp48_io_in_b = io_in_b; // @[core.scala 22:19]
endmodule
module Calc6x6(
  input         clock,
  input         reset,
  input  [15:0] io_input_mat_0,
  input  [15:0] io_input_mat_1,
  input  [15:0] io_input_mat_2,
  input  [15:0] io_input_mat_3,
  input  [15:0] io_input_mat_4,
  input  [15:0] io_input_mat_5,
  input  [15:0] io_input_mat_6,
  input  [15:0] io_input_mat_7,
  input  [15:0] io_input_mat_8,
  input  [15:0] io_input_mat_9,
  input  [15:0] io_input_mat_10,
  input  [15:0] io_input_mat_11,
  input  [15:0] io_input_mat_12,
  input  [15:0] io_input_mat_13,
  input  [15:0] io_input_mat_14,
  input  [15:0] io_input_mat_15,
  input  [15:0] io_input_mat_16,
  input  [15:0] io_input_mat_17,
  input  [15:0] io_input_mat_18,
  input  [15:0] io_input_mat_19,
  input  [15:0] io_input_mat_20,
  input  [15:0] io_input_mat_21,
  input  [15:0] io_input_mat_22,
  input  [15:0] io_input_mat_23,
  input  [15:0] io_input_mat_24,
  input  [15:0] io_input_mat_25,
  input  [15:0] io_input_mat_26,
  input  [15:0] io_input_mat_27,
  input  [15:0] io_input_mat_28,
  input  [15:0] io_input_mat_29,
  input  [15:0] io_input_mat_30,
  input  [15:0] io_input_mat_31,
  input  [15:0] io_input_mat_32,
  input  [15:0] io_input_mat_33,
  input  [15:0] io_input_mat_34,
  input  [15:0] io_input_mat_35,
  input  [1:0]  io_flag,
  input  [17:0] io_weight_real_0,
  input  [17:0] io_weight_real_1,
  input  [17:0] io_weight_real_2,
  input  [17:0] io_weight_real_3,
  input  [17:0] io_weight_real_4,
  input  [17:0] io_weight_real_5,
  input  [17:0] io_weight_real_6,
  input  [17:0] io_weight_real_7,
  input  [17:0] io_weight_real_8,
  input  [17:0] io_weight_real_9,
  input  [17:0] io_weight_real_10,
  input  [17:0] io_weight_real_11,
  input  [17:0] io_weight_real_12,
  input  [17:0] io_weight_real_13,
  input  [17:0] io_weight_real_14,
  input  [17:0] io_weight_real_15,
  input  [17:0] io_weight_comp1_0,
  input  [17:0] io_weight_comp1_1,
  input  [17:0] io_weight_comp1_2,
  input  [17:0] io_weight_comp1_3,
  input  [17:0] io_weight_comp1_4,
  input  [17:0] io_weight_comp1_5,
  input  [17:0] io_weight_comp1_6,
  input  [17:0] io_weight_comp1_7,
  input  [17:0] io_weight_comp1_8,
  input  [17:0] io_weight_comp1_9,
  input  [17:0] io_weight_comp2_0,
  input  [17:0] io_weight_comp2_1,
  input  [17:0] io_weight_comp2_2,
  input  [17:0] io_weight_comp2_3,
  input  [17:0] io_weight_comp2_4,
  input  [17:0] io_weight_comp2_5,
  input  [17:0] io_weight_comp2_6,
  input  [17:0] io_weight_comp2_7,
  input  [17:0] io_weight_comp2_8,
  input  [17:0] io_weight_comp2_9,
  input  [17:0] io_weight_comp3_0,
  input  [17:0] io_weight_comp3_1,
  input  [17:0] io_weight_comp3_2,
  input  [17:0] io_weight_comp3_3,
  input  [17:0] io_weight_comp3_4,
  input  [17:0] io_weight_comp3_5,
  input  [17:0] io_weight_comp3_6,
  input  [17:0] io_weight_comp3_7,
  input  [17:0] io_weight_comp3_8,
  input  [17:0] io_weight_comp3_9,
  output [36:0] io_output_mat_0,
  output [36:0] io_output_mat_1,
  output [36:0] io_output_mat_2,
  output [36:0] io_output_mat_3,
  output [36:0] io_output_mat_4,
  output [36:0] io_output_mat_5,
  output [36:0] io_output_mat_6,
  output [36:0] io_output_mat_7,
  output [36:0] io_output_mat_8,
  output [36:0] io_output_mat_9,
  output [36:0] io_output_mat_10,
  output [36:0] io_output_mat_11,
  output [36:0] io_output_mat_12,
  output [36:0] io_output_mat_13,
  output [36:0] io_output_mat_14,
  output [36:0] io_output_mat_15,
  input         io_valid_in,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
`endif // RANDOMIZE_REG_INIT
  wire [17:0] Core_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_1_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_1_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_1_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_1_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_2_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_2_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_2_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_2_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_3_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_3_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_3_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_3_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_4_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_4_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_4_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_4_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_5_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_5_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_5_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_5_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_6_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_6_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_6_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_6_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_7_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_7_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_7_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_7_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_8_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_8_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_8_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_8_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_9_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_9_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_9_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_9_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_10_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_10_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_10_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_10_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_11_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_11_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_11_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_11_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_12_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_12_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_12_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_12_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_13_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_13_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_13_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_13_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_14_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_14_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_14_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_14_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_15_io_w_a; // @[calc6x6.scala 64:43]
  wire [24:0] Core_15_io_in_b; // @[calc6x6.scala 64:43]
  wire  Core_15_io_flag; // @[calc6x6.scala 64:43]
  wire [42:0] Core_15_io_result; // @[calc6x6.scala 64:43]
  wire [17:0] Core_16_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_16_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_16_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_16_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_17_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_17_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_17_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_17_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_18_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_18_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_18_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_18_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_19_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_19_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_19_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_19_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_20_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_20_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_20_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_20_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_21_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_21_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_21_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_21_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_22_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_22_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_22_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_22_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_23_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_23_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_23_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_23_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_24_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_24_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_24_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_24_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_25_io_w_a; // @[calc6x6.scala 71:44]
  wire [24:0] Core_25_io_in_b; // @[calc6x6.scala 71:44]
  wire  Core_25_io_flag; // @[calc6x6.scala 71:44]
  wire [42:0] Core_25_io_result; // @[calc6x6.scala 71:44]
  wire [17:0] Core_26_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_26_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_26_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_26_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_27_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_27_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_27_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_27_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_28_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_28_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_28_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_28_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_29_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_29_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_29_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_29_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_30_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_30_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_30_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_30_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_31_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_31_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_31_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_31_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_32_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_32_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_32_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_32_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_33_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_33_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_33_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_33_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_34_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_34_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_34_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_34_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_35_io_w_a; // @[calc6x6.scala 72:44]
  wire [24:0] Core_35_io_in_b; // @[calc6x6.scala 72:44]
  wire  Core_35_io_flag; // @[calc6x6.scala 72:44]
  wire [42:0] Core_35_io_result; // @[calc6x6.scala 72:44]
  wire [17:0] Core_36_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_36_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_36_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_36_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_37_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_37_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_37_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_37_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_38_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_38_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_38_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_38_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_39_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_39_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_39_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_39_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_40_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_40_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_40_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_40_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_41_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_41_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_41_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_41_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_42_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_42_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_42_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_42_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_43_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_43_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_43_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_43_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_44_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_44_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_44_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_44_io_result; // @[calc6x6.scala 73:44]
  wire [17:0] Core_45_io_w_a; // @[calc6x6.scala 73:44]
  wire [24:0] Core_45_io_in_b; // @[calc6x6.scala 73:44]
  wire  Core_45_io_flag; // @[calc6x6.scala 73:44]
  wire [42:0] Core_45_io_result; // @[calc6x6.scala 73:44]
  reg [17:0] reg1_mat_real_0; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_1; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_2; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_3; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_4; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_5; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_6; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_7; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_8; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_9; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_10; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_11; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_12; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_13; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_14; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_15; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_16; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_17; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_18; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_19; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_20; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_21; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_22; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_23; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_30; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_31; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_32; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_33; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_34; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_real_35; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_comp_0; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_comp_1; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_comp_2; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_comp_3; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_comp_4; // @[calc6x6.scala 91:23]
  reg [17:0] reg1_mat_comp_5; // @[calc6x6.scala 91:23]
  reg [19:0] reg2_mat_real_0; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_1; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_2; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_3; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_5; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_6; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_7; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_8; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_9; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_11; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_12; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_13; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_14; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_15; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_17; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_18; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_19; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_20; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_21; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_22; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_23; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_30; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_31; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_32; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_33; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_real_35; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_0; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_1; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_2; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_3; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_4; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_5; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_6; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_7; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_8; // @[calc6x6.scala 92:23]
  reg [19:0] reg2_mat_comp_9; // @[calc6x6.scala 92:23]
  reg [37:0] w3_mat_real_0; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_1; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_2; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_3; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_4; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_5; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_6; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_7; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_8; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_9; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_10; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_11; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_12; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_13; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_14; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_15; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_16; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_17; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_18; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_19; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_20; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_21; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_22; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_23; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_24; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_25; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_26; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_27; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_28; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_29; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_30; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_31; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_32; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_33; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_34; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_real_35; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_3; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_4; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_9; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_10; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_15; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_16; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_18; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_19; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_20; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_21; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_22; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_23; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_24; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_25; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_26; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_27; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_28; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_29; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_33; // @[calc6x6.scala 93:21]
  reg [37:0] w3_mat_comp_34; // @[calc6x6.scala 93:21]
  reg [37:0] reg3_mat_real_0; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_1; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_2; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_3; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_4; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_5; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_6; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_7; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_8; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_9; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_10; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_11; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_12; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_13; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_14; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_15; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_16; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_17; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_18; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_19; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_20; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_21; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_22; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_real_23; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_comp_3; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_comp_4; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_comp_9; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_comp_10; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_comp_15; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_comp_16; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_comp_21; // @[calc6x6.scala 94:23]
  reg [37:0] reg3_mat_comp_22; // @[calc6x6.scala 94:23]
  reg  valid_reg_0; // @[calc6x6.scala 172:28]
  reg  valid_reg_1; // @[calc6x6.scala 172:28]
  reg  valid_reg_2; // @[calc6x6.scala 172:28]
  reg  valid_reg_3; // @[calc6x6.scala 172:28]
  wire [16:0] _reg1_mat_real_0_T = $signed(io_input_mat_0) - $signed(io_input_mat_24); // @[calc6x6.scala 110:56]
  wire [16:0] _reg1_mat_real_6_T = $signed(io_input_mat_6) + $signed(io_input_mat_12); // @[calc6x6.scala 111:56]
  wire [16:0] _GEN_632 = {{1{io_input_mat_18[15]}},io_input_mat_18}; // @[calc6x6.scala 111:74]
  wire [17:0] _reg1_mat_real_6_T_1 = $signed(_reg1_mat_real_6_T) + $signed(_GEN_632); // @[calc6x6.scala 111:74]
  wire [17:0] _GEN_633 = {{2{io_input_mat_24[15]}},io_input_mat_24}; // @[calc6x6.scala 111:92]
  wire [18:0] _reg1_mat_real_6_T_2 = $signed(_reg1_mat_real_6_T_1) + $signed(_GEN_633); // @[calc6x6.scala 111:92]
  wire [15:0] _reg1_mat_real_12_T_2 = 16'sh0 - $signed(io_input_mat_6); // @[calc6x6.scala 112:40]
  wire [16:0] _reg1_mat_real_12_T_3 = $signed(_reg1_mat_real_12_T_2) + $signed(io_input_mat_12); // @[calc6x6.scala 112:57]
  wire [17:0] _reg1_mat_real_12_T_4 = $signed(_reg1_mat_real_12_T_3) - $signed(_GEN_632); // @[calc6x6.scala 112:75]
  wire [18:0] _reg1_mat_real_12_T_5 = $signed(_reg1_mat_real_12_T_4) + $signed(_GEN_633); // @[calc6x6.scala 112:93]
  wire [15:0] _reg1_mat_real_18_T_2 = 16'sh0 - $signed(io_input_mat_12); // @[calc6x6.scala 113:40]
  wire [16:0] _reg1_mat_real_18_T_3 = $signed(_reg1_mat_real_18_T_2) + $signed(io_input_mat_24); // @[calc6x6.scala 113:57]
  wire [16:0] _reg1_mat_real_30_T_3 = $signed(_reg1_mat_real_12_T_2) + $signed(io_input_mat_30); // @[calc6x6.scala 115:57]
  wire [16:0] _reg1_mat_comp_0_T_3 = $signed(_reg1_mat_real_12_T_2) + $signed(io_input_mat_18); // @[calc6x6.scala 117:57]
  wire [16:0] _reg1_mat_real_1_T = $signed(io_input_mat_1) - $signed(io_input_mat_25); // @[calc6x6.scala 110:56]
  wire [16:0] _reg1_mat_real_7_T = $signed(io_input_mat_7) + $signed(io_input_mat_13); // @[calc6x6.scala 111:56]
  wire [16:0] _GEN_636 = {{1{io_input_mat_19[15]}},io_input_mat_19}; // @[calc6x6.scala 111:74]
  wire [17:0] _reg1_mat_real_7_T_1 = $signed(_reg1_mat_real_7_T) + $signed(_GEN_636); // @[calc6x6.scala 111:74]
  wire [17:0] _GEN_637 = {{2{io_input_mat_25[15]}},io_input_mat_25}; // @[calc6x6.scala 111:92]
  wire [18:0] _reg1_mat_real_7_T_2 = $signed(_reg1_mat_real_7_T_1) + $signed(_GEN_637); // @[calc6x6.scala 111:92]
  wire [15:0] _reg1_mat_real_13_T_2 = 16'sh0 - $signed(io_input_mat_7); // @[calc6x6.scala 112:40]
  wire [16:0] _reg1_mat_real_13_T_3 = $signed(_reg1_mat_real_13_T_2) + $signed(io_input_mat_13); // @[calc6x6.scala 112:57]
  wire [17:0] _reg1_mat_real_13_T_4 = $signed(_reg1_mat_real_13_T_3) - $signed(_GEN_636); // @[calc6x6.scala 112:75]
  wire [18:0] _reg1_mat_real_13_T_5 = $signed(_reg1_mat_real_13_T_4) + $signed(_GEN_637); // @[calc6x6.scala 112:93]
  wire [15:0] _reg1_mat_real_19_T_2 = 16'sh0 - $signed(io_input_mat_13); // @[calc6x6.scala 113:40]
  wire [16:0] _reg1_mat_real_19_T_3 = $signed(_reg1_mat_real_19_T_2) + $signed(io_input_mat_25); // @[calc6x6.scala 113:57]
  wire [16:0] _reg1_mat_real_31_T_3 = $signed(_reg1_mat_real_13_T_2) + $signed(io_input_mat_31); // @[calc6x6.scala 115:57]
  wire [16:0] _reg1_mat_comp_1_T_3 = $signed(_reg1_mat_real_13_T_2) + $signed(io_input_mat_19); // @[calc6x6.scala 117:57]
  wire [16:0] _reg1_mat_real_2_T = $signed(io_input_mat_2) - $signed(io_input_mat_26); // @[calc6x6.scala 110:56]
  wire [16:0] _reg1_mat_real_8_T = $signed(io_input_mat_8) + $signed(io_input_mat_14); // @[calc6x6.scala 111:56]
  wire [16:0] _GEN_640 = {{1{io_input_mat_20[15]}},io_input_mat_20}; // @[calc6x6.scala 111:74]
  wire [17:0] _reg1_mat_real_8_T_1 = $signed(_reg1_mat_real_8_T) + $signed(_GEN_640); // @[calc6x6.scala 111:74]
  wire [17:0] _GEN_641 = {{2{io_input_mat_26[15]}},io_input_mat_26}; // @[calc6x6.scala 111:92]
  wire [18:0] _reg1_mat_real_8_T_2 = $signed(_reg1_mat_real_8_T_1) + $signed(_GEN_641); // @[calc6x6.scala 111:92]
  wire [15:0] _reg1_mat_real_14_T_2 = 16'sh0 - $signed(io_input_mat_8); // @[calc6x6.scala 112:40]
  wire [16:0] _reg1_mat_real_14_T_3 = $signed(_reg1_mat_real_14_T_2) + $signed(io_input_mat_14); // @[calc6x6.scala 112:57]
  wire [17:0] _reg1_mat_real_14_T_4 = $signed(_reg1_mat_real_14_T_3) - $signed(_GEN_640); // @[calc6x6.scala 112:75]
  wire [18:0] _reg1_mat_real_14_T_5 = $signed(_reg1_mat_real_14_T_4) + $signed(_GEN_641); // @[calc6x6.scala 112:93]
  wire [15:0] _reg1_mat_real_20_T_2 = 16'sh0 - $signed(io_input_mat_14); // @[calc6x6.scala 113:40]
  wire [16:0] _reg1_mat_real_20_T_3 = $signed(_reg1_mat_real_20_T_2) + $signed(io_input_mat_26); // @[calc6x6.scala 113:57]
  wire [16:0] _reg1_mat_real_32_T_3 = $signed(_reg1_mat_real_14_T_2) + $signed(io_input_mat_32); // @[calc6x6.scala 115:57]
  wire [16:0] _reg1_mat_comp_2_T_3 = $signed(_reg1_mat_real_14_T_2) + $signed(io_input_mat_20); // @[calc6x6.scala 117:57]
  wire [16:0] _reg1_mat_real_3_T = $signed(io_input_mat_3) - $signed(io_input_mat_27); // @[calc6x6.scala 110:56]
  wire [16:0] _reg1_mat_real_9_T = $signed(io_input_mat_9) + $signed(io_input_mat_15); // @[calc6x6.scala 111:56]
  wire [16:0] _GEN_644 = {{1{io_input_mat_21[15]}},io_input_mat_21}; // @[calc6x6.scala 111:74]
  wire [17:0] _reg1_mat_real_9_T_1 = $signed(_reg1_mat_real_9_T) + $signed(_GEN_644); // @[calc6x6.scala 111:74]
  wire [17:0] _GEN_645 = {{2{io_input_mat_27[15]}},io_input_mat_27}; // @[calc6x6.scala 111:92]
  wire [18:0] _reg1_mat_real_9_T_2 = $signed(_reg1_mat_real_9_T_1) + $signed(_GEN_645); // @[calc6x6.scala 111:92]
  wire [15:0] _reg1_mat_real_15_T_2 = 16'sh0 - $signed(io_input_mat_9); // @[calc6x6.scala 112:40]
  wire [16:0] _reg1_mat_real_15_T_3 = $signed(_reg1_mat_real_15_T_2) + $signed(io_input_mat_15); // @[calc6x6.scala 112:57]
  wire [17:0] _reg1_mat_real_15_T_4 = $signed(_reg1_mat_real_15_T_3) - $signed(_GEN_644); // @[calc6x6.scala 112:75]
  wire [18:0] _reg1_mat_real_15_T_5 = $signed(_reg1_mat_real_15_T_4) + $signed(_GEN_645); // @[calc6x6.scala 112:93]
  wire [15:0] _reg1_mat_real_21_T_2 = 16'sh0 - $signed(io_input_mat_15); // @[calc6x6.scala 113:40]
  wire [16:0] _reg1_mat_real_21_T_3 = $signed(_reg1_mat_real_21_T_2) + $signed(io_input_mat_27); // @[calc6x6.scala 113:57]
  wire [16:0] _reg1_mat_real_33_T_3 = $signed(_reg1_mat_real_15_T_2) + $signed(io_input_mat_33); // @[calc6x6.scala 115:57]
  wire [16:0] _reg1_mat_comp_3_T_3 = $signed(_reg1_mat_real_15_T_2) + $signed(io_input_mat_21); // @[calc6x6.scala 117:57]
  wire [16:0] _reg1_mat_real_4_T = $signed(io_input_mat_4) - $signed(io_input_mat_28); // @[calc6x6.scala 110:56]
  wire [16:0] _reg1_mat_real_10_T = $signed(io_input_mat_10) + $signed(io_input_mat_16); // @[calc6x6.scala 111:56]
  wire [16:0] _GEN_648 = {{1{io_input_mat_22[15]}},io_input_mat_22}; // @[calc6x6.scala 111:74]
  wire [17:0] _reg1_mat_real_10_T_1 = $signed(_reg1_mat_real_10_T) + $signed(_GEN_648); // @[calc6x6.scala 111:74]
  wire [17:0] _GEN_649 = {{2{io_input_mat_28[15]}},io_input_mat_28}; // @[calc6x6.scala 111:92]
  wire [18:0] _reg1_mat_real_10_T_2 = $signed(_reg1_mat_real_10_T_1) + $signed(_GEN_649); // @[calc6x6.scala 111:92]
  wire [15:0] _reg1_mat_real_16_T_2 = 16'sh0 - $signed(io_input_mat_10); // @[calc6x6.scala 112:40]
  wire [16:0] _reg1_mat_real_16_T_3 = $signed(_reg1_mat_real_16_T_2) + $signed(io_input_mat_16); // @[calc6x6.scala 112:57]
  wire [17:0] _reg1_mat_real_16_T_4 = $signed(_reg1_mat_real_16_T_3) - $signed(_GEN_648); // @[calc6x6.scala 112:75]
  wire [18:0] _reg1_mat_real_16_T_5 = $signed(_reg1_mat_real_16_T_4) + $signed(_GEN_649); // @[calc6x6.scala 112:93]
  wire [15:0] _reg1_mat_real_22_T_2 = 16'sh0 - $signed(io_input_mat_16); // @[calc6x6.scala 113:40]
  wire [16:0] _reg1_mat_real_22_T_3 = $signed(_reg1_mat_real_22_T_2) + $signed(io_input_mat_28); // @[calc6x6.scala 113:57]
  wire [16:0] _reg1_mat_real_34_T_3 = $signed(_reg1_mat_real_16_T_2) + $signed(io_input_mat_34); // @[calc6x6.scala 115:57]
  wire [16:0] _reg1_mat_comp_4_T_3 = $signed(_reg1_mat_real_16_T_2) + $signed(io_input_mat_22); // @[calc6x6.scala 117:57]
  wire [16:0] _reg1_mat_real_5_T = $signed(io_input_mat_5) - $signed(io_input_mat_29); // @[calc6x6.scala 110:56]
  wire [16:0] _reg1_mat_real_11_T = $signed(io_input_mat_11) + $signed(io_input_mat_17); // @[calc6x6.scala 111:56]
  wire [16:0] _GEN_652 = {{1{io_input_mat_23[15]}},io_input_mat_23}; // @[calc6x6.scala 111:74]
  wire [17:0] _reg1_mat_real_11_T_1 = $signed(_reg1_mat_real_11_T) + $signed(_GEN_652); // @[calc6x6.scala 111:74]
  wire [17:0] _GEN_653 = {{2{io_input_mat_29[15]}},io_input_mat_29}; // @[calc6x6.scala 111:92]
  wire [18:0] _reg1_mat_real_11_T_2 = $signed(_reg1_mat_real_11_T_1) + $signed(_GEN_653); // @[calc6x6.scala 111:92]
  wire [15:0] _reg1_mat_real_17_T_2 = 16'sh0 - $signed(io_input_mat_11); // @[calc6x6.scala 112:40]
  wire [16:0] _reg1_mat_real_17_T_3 = $signed(_reg1_mat_real_17_T_2) + $signed(io_input_mat_17); // @[calc6x6.scala 112:57]
  wire [17:0] _reg1_mat_real_17_T_4 = $signed(_reg1_mat_real_17_T_3) - $signed(_GEN_652); // @[calc6x6.scala 112:75]
  wire [18:0] _reg1_mat_real_17_T_5 = $signed(_reg1_mat_real_17_T_4) + $signed(_GEN_653); // @[calc6x6.scala 112:93]
  wire [15:0] _reg1_mat_real_23_T_2 = 16'sh0 - $signed(io_input_mat_17); // @[calc6x6.scala 113:40]
  wire [16:0] _reg1_mat_real_23_T_3 = $signed(_reg1_mat_real_23_T_2) + $signed(io_input_mat_29); // @[calc6x6.scala 113:57]
  wire [16:0] _reg1_mat_real_35_T_3 = $signed(_reg1_mat_real_17_T_2) + $signed(io_input_mat_35); // @[calc6x6.scala 115:57]
  wire [16:0] _reg1_mat_comp_5_T_3 = $signed(_reg1_mat_real_17_T_2) + $signed(io_input_mat_23); // @[calc6x6.scala 117:57]
  wire [18:0] _reg2_mat_real_0_T = $signed(reg1_mat_real_0) - $signed(reg1_mat_real_4); // @[calc6x6.scala 124:61]
  wire [18:0] _reg2_mat_real_1_T = $signed(reg1_mat_real_1) + $signed(reg1_mat_real_2); // @[calc6x6.scala 125:61]
  wire [18:0] _GEN_656 = {{1{reg1_mat_real_3[17]}},reg1_mat_real_3}; // @[calc6x6.scala 125:84]
  wire [19:0] _reg2_mat_real_1_T_1 = $signed(_reg2_mat_real_1_T) + $signed(_GEN_656); // @[calc6x6.scala 125:84]
  wire [19:0] _GEN_657 = {{2{reg1_mat_real_4[17]}},reg1_mat_real_4}; // @[calc6x6.scala 125:107]
  wire [20:0] _reg2_mat_real_1_T_2 = $signed(_reg2_mat_real_1_T_1) + $signed(_GEN_657); // @[calc6x6.scala 125:107]
  wire [17:0] _reg2_mat_real_2_T_2 = 18'sh0 - $signed(reg1_mat_real_1); // @[calc6x6.scala 126:40]
  wire [18:0] _reg2_mat_real_2_T_3 = $signed(_reg2_mat_real_2_T_2) + $signed(reg1_mat_real_2); // @[calc6x6.scala 126:62]
  wire [19:0] _reg2_mat_real_2_T_4 = $signed(_reg2_mat_real_2_T_3) - $signed(_GEN_656); // @[calc6x6.scala 126:85]
  wire [20:0] _reg2_mat_real_2_T_5 = $signed(_reg2_mat_real_2_T_4) + $signed(_GEN_657); // @[calc6x6.scala 126:108]
  wire [17:0] _reg2_mat_real_3_T_2 = 18'sh0 - $signed(reg1_mat_real_2); // @[calc6x6.scala 127:158]
  wire [18:0] _reg2_mat_real_3_T_3 = $signed(_reg2_mat_real_3_T_2) + $signed(reg1_mat_real_4); // @[calc6x6.scala 127:180]
  wire [18:0] _reg2_mat_real_5_T_3 = $signed(_reg2_mat_real_2_T_2) + $signed(reg1_mat_real_5); // @[calc6x6.scala 129:62]
  wire [18:0] _reg2_mat_real_6_T = $signed(reg1_mat_real_6) - $signed(reg1_mat_real_10); // @[calc6x6.scala 124:61]
  wire [18:0] _reg2_mat_real_7_T = $signed(reg1_mat_real_7) + $signed(reg1_mat_real_8); // @[calc6x6.scala 125:61]
  wire [18:0] _GEN_660 = {{1{reg1_mat_real_9[17]}},reg1_mat_real_9}; // @[calc6x6.scala 125:84]
  wire [19:0] _reg2_mat_real_7_T_1 = $signed(_reg2_mat_real_7_T) + $signed(_GEN_660); // @[calc6x6.scala 125:84]
  wire [19:0] _GEN_661 = {{2{reg1_mat_real_10[17]}},reg1_mat_real_10}; // @[calc6x6.scala 125:107]
  wire [20:0] _reg2_mat_real_7_T_2 = $signed(_reg2_mat_real_7_T_1) + $signed(_GEN_661); // @[calc6x6.scala 125:107]
  wire [17:0] _reg2_mat_real_8_T_2 = 18'sh0 - $signed(reg1_mat_real_7); // @[calc6x6.scala 126:40]
  wire [18:0] _reg2_mat_real_8_T_3 = $signed(_reg2_mat_real_8_T_2) + $signed(reg1_mat_real_8); // @[calc6x6.scala 126:62]
  wire [19:0] _reg2_mat_real_8_T_4 = $signed(_reg2_mat_real_8_T_3) - $signed(_GEN_660); // @[calc6x6.scala 126:85]
  wire [20:0] _reg2_mat_real_8_T_5 = $signed(_reg2_mat_real_8_T_4) + $signed(_GEN_661); // @[calc6x6.scala 126:108]
  wire [17:0] _reg2_mat_real_9_T_2 = 18'sh0 - $signed(reg1_mat_real_8); // @[calc6x6.scala 127:158]
  wire [18:0] _reg2_mat_real_9_T_3 = $signed(_reg2_mat_real_9_T_2) + $signed(reg1_mat_real_10); // @[calc6x6.scala 127:180]
  wire [18:0] _reg2_mat_real_11_T_3 = $signed(_reg2_mat_real_8_T_2) + $signed(reg1_mat_real_11); // @[calc6x6.scala 129:62]
  wire [18:0] _reg2_mat_real_12_T = $signed(reg1_mat_real_12) - $signed(reg1_mat_real_16); // @[calc6x6.scala 124:61]
  wire [18:0] _reg2_mat_real_13_T = $signed(reg1_mat_real_13) + $signed(reg1_mat_real_14); // @[calc6x6.scala 125:61]
  wire [18:0] _GEN_664 = {{1{reg1_mat_real_15[17]}},reg1_mat_real_15}; // @[calc6x6.scala 125:84]
  wire [19:0] _reg2_mat_real_13_T_1 = $signed(_reg2_mat_real_13_T) + $signed(_GEN_664); // @[calc6x6.scala 125:84]
  wire [19:0] _GEN_665 = {{2{reg1_mat_real_16[17]}},reg1_mat_real_16}; // @[calc6x6.scala 125:107]
  wire [20:0] _reg2_mat_real_13_T_2 = $signed(_reg2_mat_real_13_T_1) + $signed(_GEN_665); // @[calc6x6.scala 125:107]
  wire [17:0] _reg2_mat_real_14_T_2 = 18'sh0 - $signed(reg1_mat_real_13); // @[calc6x6.scala 126:40]
  wire [18:0] _reg2_mat_real_14_T_3 = $signed(_reg2_mat_real_14_T_2) + $signed(reg1_mat_real_14); // @[calc6x6.scala 126:62]
  wire [19:0] _reg2_mat_real_14_T_4 = $signed(_reg2_mat_real_14_T_3) - $signed(_GEN_664); // @[calc6x6.scala 126:85]
  wire [20:0] _reg2_mat_real_14_T_5 = $signed(_reg2_mat_real_14_T_4) + $signed(_GEN_665); // @[calc6x6.scala 126:108]
  wire [17:0] _reg2_mat_real_15_T_2 = 18'sh0 - $signed(reg1_mat_real_14); // @[calc6x6.scala 127:158]
  wire [18:0] _reg2_mat_real_15_T_3 = $signed(_reg2_mat_real_15_T_2) + $signed(reg1_mat_real_16); // @[calc6x6.scala 127:180]
  wire [18:0] _reg2_mat_real_17_T_3 = $signed(_reg2_mat_real_14_T_2) + $signed(reg1_mat_real_17); // @[calc6x6.scala 129:62]
  wire [18:0] _reg2_mat_real_18_T = $signed(reg1_mat_real_18) - $signed(reg1_mat_real_22); // @[calc6x6.scala 124:61]
  wire [18:0] _reg2_mat_real_19_T = $signed(reg1_mat_real_19) + $signed(reg1_mat_real_20); // @[calc6x6.scala 125:61]
  wire [18:0] _GEN_668 = {{1{reg1_mat_real_21[17]}},reg1_mat_real_21}; // @[calc6x6.scala 125:84]
  wire [19:0] _reg2_mat_real_19_T_1 = $signed(_reg2_mat_real_19_T) + $signed(_GEN_668); // @[calc6x6.scala 125:84]
  wire [19:0] _GEN_669 = {{2{reg1_mat_real_22[17]}},reg1_mat_real_22}; // @[calc6x6.scala 125:107]
  wire [20:0] _reg2_mat_real_19_T_2 = $signed(_reg2_mat_real_19_T_1) + $signed(_GEN_669); // @[calc6x6.scala 125:107]
  wire [17:0] _reg2_mat_real_20_T_2 = 18'sh0 - $signed(reg1_mat_real_19); // @[calc6x6.scala 126:40]
  wire [18:0] _reg2_mat_real_20_T_3 = $signed(_reg2_mat_real_20_T_2) + $signed(reg1_mat_real_20); // @[calc6x6.scala 126:62]
  wire [19:0] _reg2_mat_real_20_T_4 = $signed(_reg2_mat_real_20_T_3) - $signed(_GEN_668); // @[calc6x6.scala 126:85]
  wire [20:0] _reg2_mat_real_20_T_5 = $signed(_reg2_mat_real_20_T_4) + $signed(_GEN_669); // @[calc6x6.scala 126:108]
  wire [17:0] _reg2_mat_real_21_T_2 = 18'sh0 - $signed(reg1_mat_real_20); // @[calc6x6.scala 127:57]
  wire [18:0] _reg2_mat_real_21_T_3 = $signed(_reg2_mat_real_21_T_2) + $signed(reg1_mat_real_22); // @[calc6x6.scala 127:79]
  wire [18:0] _GEN_672 = {{1{reg1_mat_comp_3[17]}},reg1_mat_comp_3}; // @[calc6x6.scala 127:102]
  wire [19:0] _reg2_mat_real_21_T_4 = $signed(_reg2_mat_real_21_T_3) - $signed(_GEN_672); // @[calc6x6.scala 127:102]
  wire [19:0] _GEN_673 = {{2{reg1_mat_comp_1[17]}},reg1_mat_comp_1}; // @[calc6x6.scala 127:127]
  wire [20:0] _reg2_mat_real_21_T_5 = $signed(_reg2_mat_real_21_T_4) + $signed(_GEN_673); // @[calc6x6.scala 127:127]
  wire [19:0] _reg2_mat_real_22_T_4 = $signed(_reg2_mat_real_21_T_3) + $signed(_GEN_672); // @[calc6x6.scala 128:102]
  wire [20:0] _reg2_mat_real_22_T_5 = $signed(_reg2_mat_real_22_T_4) - $signed(_GEN_673); // @[calc6x6.scala 128:127]
  wire [18:0] _reg2_mat_real_23_T_3 = $signed(_reg2_mat_real_20_T_2) + $signed(reg1_mat_real_23); // @[calc6x6.scala 129:62]
  wire [18:0] _reg2_mat_real_30_T = $signed(reg1_mat_real_30) - $signed(reg1_mat_real_34); // @[calc6x6.scala 124:61]
  wire [18:0] _reg2_mat_real_31_T = $signed(reg1_mat_real_31) + $signed(reg1_mat_real_32); // @[calc6x6.scala 125:61]
  wire [18:0] _GEN_684 = {{1{reg1_mat_real_33[17]}},reg1_mat_real_33}; // @[calc6x6.scala 125:84]
  wire [19:0] _reg2_mat_real_31_T_1 = $signed(_reg2_mat_real_31_T) + $signed(_GEN_684); // @[calc6x6.scala 125:84]
  wire [19:0] _GEN_685 = {{2{reg1_mat_real_34[17]}},reg1_mat_real_34}; // @[calc6x6.scala 125:107]
  wire [20:0] _reg2_mat_real_31_T_2 = $signed(_reg2_mat_real_31_T_1) + $signed(_GEN_685); // @[calc6x6.scala 125:107]
  wire [17:0] _reg2_mat_real_32_T_2 = 18'sh0 - $signed(reg1_mat_real_31); // @[calc6x6.scala 126:40]
  wire [18:0] _reg2_mat_real_32_T_3 = $signed(_reg2_mat_real_32_T_2) + $signed(reg1_mat_real_32); // @[calc6x6.scala 126:62]
  wire [19:0] _reg2_mat_real_32_T_4 = $signed(_reg2_mat_real_32_T_3) - $signed(_GEN_684); // @[calc6x6.scala 126:85]
  wire [20:0] _reg2_mat_real_32_T_5 = $signed(_reg2_mat_real_32_T_4) + $signed(_GEN_685); // @[calc6x6.scala 126:108]
  wire [17:0] _reg2_mat_real_33_T_2 = 18'sh0 - $signed(reg1_mat_real_32); // @[calc6x6.scala 127:158]
  wire [18:0] _reg2_mat_real_33_T_3 = $signed(_reg2_mat_real_33_T_2) + $signed(reg1_mat_real_34); // @[calc6x6.scala 127:180]
  wire [18:0] _reg2_mat_real_35_T_3 = $signed(_reg2_mat_real_32_T_2) + $signed(reg1_mat_real_35); // @[calc6x6.scala 129:62]
  wire [18:0] _reg2_mat_comp_0_T = $signed(reg1_mat_comp_0) - $signed(reg1_mat_comp_4); // @[calc6x6.scala 132:50]
  wire [18:0] _reg2_mat_comp_1_T = $signed(reg1_mat_comp_1) + $signed(reg1_mat_comp_2); // @[calc6x6.scala 133:50]
  wire [19:0] _reg2_mat_comp_1_T_1 = $signed(_reg2_mat_comp_1_T) + $signed(_GEN_672); // @[calc6x6.scala 133:73]
  wire [19:0] _GEN_689 = {{2{reg1_mat_comp_4[17]}},reg1_mat_comp_4}; // @[calc6x6.scala 133:96]
  wire [20:0] _reg2_mat_comp_1_T_2 = $signed(_reg2_mat_comp_1_T_1) + $signed(_GEN_689); // @[calc6x6.scala 133:96]
  wire [17:0] _reg2_mat_comp_2_T_2 = 18'sh0 - $signed(reg1_mat_comp_1); // @[calc6x6.scala 134:29]
  wire [18:0] _reg2_mat_comp_2_T_3 = $signed(_reg2_mat_comp_2_T_2) + $signed(reg1_mat_comp_2); // @[calc6x6.scala 134:51]
  wire [19:0] _reg2_mat_comp_2_T_4 = $signed(_reg2_mat_comp_2_T_3) - $signed(_GEN_672); // @[calc6x6.scala 134:74]
  wire [20:0] _reg2_mat_comp_2_T_5 = $signed(_reg2_mat_comp_2_T_4) + $signed(_GEN_689); // @[calc6x6.scala 134:97]
  wire [17:0] _reg2_mat_comp_3_T_2 = 18'sh0 - $signed(reg1_mat_comp_2); // @[calc6x6.scala 135:29]
  wire [18:0] _reg2_mat_comp_3_T_3 = $signed(_reg2_mat_comp_3_T_2) + $signed(reg1_mat_comp_4); // @[calc6x6.scala 135:51]
  wire [18:0] _GEN_692 = {{1{reg1_mat_real_19[17]}},reg1_mat_real_19}; // @[calc6x6.scala 135:74]
  wire [19:0] _reg2_mat_comp_3_T_4 = $signed(_reg2_mat_comp_3_T_3) - $signed(_GEN_692); // @[calc6x6.scala 135:74]
  wire [19:0] _GEN_693 = {{2{reg1_mat_real_21[17]}},reg1_mat_real_21}; // @[calc6x6.scala 135:97]
  wire [20:0] _reg2_mat_comp_3_T_5 = $signed(_reg2_mat_comp_3_T_4) + $signed(_GEN_693); // @[calc6x6.scala 135:97]
  wire [19:0] _reg2_mat_comp_4_T_4 = $signed(_reg2_mat_comp_3_T_3) + $signed(_GEN_692); // @[calc6x6.scala 136:74]
  wire [20:0] _reg2_mat_comp_4_T_5 = $signed(_reg2_mat_comp_4_T_4) - $signed(_GEN_693); // @[calc6x6.scala 136:97]
  wire [18:0] _reg2_mat_comp_5_T_3 = $signed(_reg2_mat_comp_2_T_2) + $signed(reg1_mat_comp_5); // @[calc6x6.scala 137:51]
  wire [18:0] _reg2_mat_comp_6_T_3 = $signed(_reg2_mat_real_2_T_2) + $signed(reg1_mat_real_3); // @[calc6x6.scala 140:51]
  wire [18:0] _reg2_mat_comp_7_T_3 = $signed(_reg2_mat_real_8_T_2) + $signed(reg1_mat_real_9); // @[calc6x6.scala 141:51]
  wire [18:0] _reg2_mat_comp_8_T_3 = $signed(_reg2_mat_real_14_T_2) + $signed(reg1_mat_real_15); // @[calc6x6.scala 142:51]
  wire [18:0] _reg2_mat_comp_9_T_3 = $signed(_reg2_mat_real_32_T_2) + $signed(reg1_mat_real_33); // @[calc6x6.scala 143:51]
  wire [37:0] _reg3_mat_real_0_T_2 = $signed(w3_mat_real_6) + $signed(w3_mat_real_12); // @[calc6x6.scala 148:85]
  wire [37:0] _reg3_mat_real_0_T_5 = $signed(_reg3_mat_real_0_T_2) + $signed(w3_mat_real_18); // @[calc6x6.scala 149:62]
  wire [37:0] _reg3_mat_real_0_T_8 = $signed(_reg3_mat_real_0_T_5) + $signed(w3_mat_real_24); // @[calc6x6.scala 149:84]
  wire [35:0] _GEN_696 = _reg3_mat_real_0_T_8[37:2]; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_0_T_9 = {{2{_GEN_696[35]}},_GEN_696}; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_0_T_12 = $signed(w3_mat_real_0) + $signed(_reg3_mat_real_0_T_9); // @[calc6x6.scala 148:61]
  wire [37:0] _reg3_mat_real_6_T_2 = $signed(w3_mat_real_6) - $signed(w3_mat_real_12); // @[calc6x6.scala 150:62]
  wire [37:0] _reg3_mat_real_6_T_5 = $signed(_reg3_mat_real_6_T_2) - $signed(w3_mat_comp_18); // @[calc6x6.scala 150:84]
  wire [37:0] _reg3_mat_real_6_T_8 = $signed(_reg3_mat_real_6_T_5) + $signed(w3_mat_comp_24); // @[calc6x6.scala 150:106]
  wire [35:0] _GEN_697 = _reg3_mat_real_6_T_8[37:2]; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_6_T_9 = {{2{_GEN_697[35]}},_GEN_697}; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_12_T_5 = $signed(_reg3_mat_real_0_T_2) - $signed(w3_mat_real_18); // @[calc6x6.scala 151:84]
  wire [37:0] _reg3_mat_real_12_T_8 = $signed(_reg3_mat_real_12_T_5) - $signed(w3_mat_real_24); // @[calc6x6.scala 151:106]
  wire [35:0] _GEN_698 = _reg3_mat_real_12_T_8[37:2]; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_12_T_9 = {{2{_GEN_698[35]}},_GEN_698}; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_18_T_5 = $signed(_reg3_mat_real_6_T_2) + $signed(w3_mat_comp_18); // @[calc6x6.scala 152:85]
  wire [37:0] _reg3_mat_real_18_T_8 = $signed(_reg3_mat_real_18_T_5) - $signed(w3_mat_comp_24); // @[calc6x6.scala 152:107]
  wire [35:0] _GEN_699 = _reg3_mat_real_18_T_8[37:2]; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_18_T_9 = {{2{_GEN_699[35]}},_GEN_699}; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_18_T_12 = $signed(_reg3_mat_real_18_T_9) + $signed(w3_mat_real_30); // @[calc6x6.scala 152:136]
  wire [37:0] _reg3_mat_real_1_T_2 = $signed(w3_mat_real_7) + $signed(w3_mat_real_13); // @[calc6x6.scala 148:85]
  wire [37:0] _reg3_mat_real_1_T_5 = $signed(_reg3_mat_real_1_T_2) + $signed(w3_mat_real_19); // @[calc6x6.scala 149:62]
  wire [37:0] _reg3_mat_real_1_T_8 = $signed(_reg3_mat_real_1_T_5) + $signed(w3_mat_real_25); // @[calc6x6.scala 149:84]
  wire [35:0] _GEN_704 = _reg3_mat_real_1_T_8[37:2]; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_1_T_9 = {{2{_GEN_704[35]}},_GEN_704}; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_1_T_12 = $signed(w3_mat_real_1) + $signed(_reg3_mat_real_1_T_9); // @[calc6x6.scala 148:61]
  wire [37:0] _reg3_mat_real_7_T_2 = $signed(w3_mat_real_7) - $signed(w3_mat_real_13); // @[calc6x6.scala 150:62]
  wire [37:0] _reg3_mat_real_7_T_5 = $signed(_reg3_mat_real_7_T_2) - $signed(w3_mat_comp_19); // @[calc6x6.scala 150:84]
  wire [37:0] _reg3_mat_real_7_T_8 = $signed(_reg3_mat_real_7_T_5) + $signed(w3_mat_comp_25); // @[calc6x6.scala 150:106]
  wire [35:0] _GEN_705 = _reg3_mat_real_7_T_8[37:2]; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_7_T_9 = {{2{_GEN_705[35]}},_GEN_705}; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_13_T_5 = $signed(_reg3_mat_real_1_T_2) - $signed(w3_mat_real_19); // @[calc6x6.scala 151:84]
  wire [37:0] _reg3_mat_real_13_T_8 = $signed(_reg3_mat_real_13_T_5) - $signed(w3_mat_real_25); // @[calc6x6.scala 151:106]
  wire [35:0] _GEN_706 = _reg3_mat_real_13_T_8[37:2]; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_13_T_9 = {{2{_GEN_706[35]}},_GEN_706}; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_19_T_5 = $signed(_reg3_mat_real_7_T_2) + $signed(w3_mat_comp_19); // @[calc6x6.scala 152:85]
  wire [37:0] _reg3_mat_real_19_T_8 = $signed(_reg3_mat_real_19_T_5) - $signed(w3_mat_comp_25); // @[calc6x6.scala 152:107]
  wire [35:0] _GEN_707 = _reg3_mat_real_19_T_8[37:2]; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_19_T_9 = {{2{_GEN_707[35]}},_GEN_707}; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_19_T_12 = $signed(_reg3_mat_real_19_T_9) + $signed(w3_mat_real_31); // @[calc6x6.scala 152:136]
  wire [37:0] _reg3_mat_real_2_T_2 = $signed(w3_mat_real_8) + $signed(w3_mat_real_14); // @[calc6x6.scala 148:85]
  wire [37:0] _reg3_mat_real_2_T_5 = $signed(_reg3_mat_real_2_T_2) + $signed(w3_mat_real_20); // @[calc6x6.scala 149:62]
  wire [37:0] _reg3_mat_real_2_T_8 = $signed(_reg3_mat_real_2_T_5) + $signed(w3_mat_real_26); // @[calc6x6.scala 149:84]
  wire [35:0] _GEN_712 = _reg3_mat_real_2_T_8[37:2]; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_2_T_9 = {{2{_GEN_712[35]}},_GEN_712}; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_2_T_12 = $signed(w3_mat_real_2) + $signed(_reg3_mat_real_2_T_9); // @[calc6x6.scala 148:61]
  wire [37:0] _reg3_mat_real_8_T_2 = $signed(w3_mat_real_8) - $signed(w3_mat_real_14); // @[calc6x6.scala 150:62]
  wire [37:0] _reg3_mat_real_8_T_5 = $signed(_reg3_mat_real_8_T_2) - $signed(w3_mat_comp_20); // @[calc6x6.scala 150:84]
  wire [37:0] _reg3_mat_real_8_T_8 = $signed(_reg3_mat_real_8_T_5) + $signed(w3_mat_comp_26); // @[calc6x6.scala 150:106]
  wire [35:0] _GEN_713 = _reg3_mat_real_8_T_8[37:2]; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_8_T_9 = {{2{_GEN_713[35]}},_GEN_713}; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_14_T_5 = $signed(_reg3_mat_real_2_T_2) - $signed(w3_mat_real_20); // @[calc6x6.scala 151:84]
  wire [37:0] _reg3_mat_real_14_T_8 = $signed(_reg3_mat_real_14_T_5) - $signed(w3_mat_real_26); // @[calc6x6.scala 151:106]
  wire [35:0] _GEN_714 = _reg3_mat_real_14_T_8[37:2]; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_14_T_9 = {{2{_GEN_714[35]}},_GEN_714}; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_20_T_5 = $signed(_reg3_mat_real_8_T_2) + $signed(w3_mat_comp_20); // @[calc6x6.scala 152:85]
  wire [37:0] _reg3_mat_real_20_T_8 = $signed(_reg3_mat_real_20_T_5) - $signed(w3_mat_comp_26); // @[calc6x6.scala 152:107]
  wire [35:0] _GEN_715 = _reg3_mat_real_20_T_8[37:2]; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_20_T_9 = {{2{_GEN_715[35]}},_GEN_715}; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_20_T_12 = $signed(_reg3_mat_real_20_T_9) + $signed(w3_mat_real_32); // @[calc6x6.scala 152:136]
  wire [37:0] _reg3_mat_real_3_T_2 = $signed(w3_mat_real_9) + $signed(w3_mat_real_15); // @[calc6x6.scala 148:85]
  wire [37:0] _reg3_mat_real_3_T_5 = $signed(_reg3_mat_real_3_T_2) + $signed(w3_mat_real_21); // @[calc6x6.scala 149:62]
  wire [37:0] _reg3_mat_real_3_T_8 = $signed(_reg3_mat_real_3_T_5) + $signed(w3_mat_real_27); // @[calc6x6.scala 149:84]
  wire [35:0] _GEN_720 = _reg3_mat_real_3_T_8[37:2]; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_3_T_9 = {{2{_GEN_720[35]}},_GEN_720}; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_3_T_12 = $signed(w3_mat_real_3) + $signed(_reg3_mat_real_3_T_9); // @[calc6x6.scala 148:61]
  wire [37:0] _reg3_mat_real_9_T_2 = $signed(w3_mat_real_9) - $signed(w3_mat_real_15); // @[calc6x6.scala 150:62]
  wire [37:0] _reg3_mat_real_9_T_5 = $signed(_reg3_mat_real_9_T_2) - $signed(w3_mat_comp_21); // @[calc6x6.scala 150:84]
  wire [37:0] _reg3_mat_real_9_T_8 = $signed(_reg3_mat_real_9_T_5) + $signed(w3_mat_comp_27); // @[calc6x6.scala 150:106]
  wire [35:0] _GEN_721 = _reg3_mat_real_9_T_8[37:2]; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_9_T_9 = {{2{_GEN_721[35]}},_GEN_721}; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_15_T_5 = $signed(_reg3_mat_real_3_T_2) - $signed(w3_mat_real_21); // @[calc6x6.scala 151:84]
  wire [37:0] _reg3_mat_real_15_T_8 = $signed(_reg3_mat_real_15_T_5) - $signed(w3_mat_real_27); // @[calc6x6.scala 151:106]
  wire [35:0] _GEN_722 = _reg3_mat_real_15_T_8[37:2]; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_15_T_9 = {{2{_GEN_722[35]}},_GEN_722}; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_21_T_5 = $signed(_reg3_mat_real_9_T_2) + $signed(w3_mat_comp_21); // @[calc6x6.scala 152:85]
  wire [37:0] _reg3_mat_real_21_T_8 = $signed(_reg3_mat_real_21_T_5) - $signed(w3_mat_comp_27); // @[calc6x6.scala 152:107]
  wire [35:0] _GEN_723 = _reg3_mat_real_21_T_8[37:2]; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_21_T_9 = {{2{_GEN_723[35]}},_GEN_723}; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_21_T_12 = $signed(_reg3_mat_real_21_T_9) + $signed(w3_mat_real_33); // @[calc6x6.scala 152:136]
  wire [37:0] _reg3_mat_comp_3_T_2 = $signed(w3_mat_comp_9) + $signed(w3_mat_comp_15); // @[calc6x6.scala 154:85]
  wire [37:0] _reg3_mat_comp_3_T_5 = $signed(_reg3_mat_comp_3_T_2) + $signed(w3_mat_comp_21); // @[calc6x6.scala 155:62]
  wire [37:0] _reg3_mat_comp_3_T_8 = $signed(_reg3_mat_comp_3_T_5) + $signed(w3_mat_comp_27); // @[calc6x6.scala 155:84]
  wire [35:0] _GEN_724 = _reg3_mat_comp_3_T_8[37:2]; // @[calc6x6.scala 155:107]
  wire [37:0] _reg3_mat_comp_3_T_9 = {{2{_GEN_724[35]}},_GEN_724}; // @[calc6x6.scala 155:107]
  wire [37:0] _reg3_mat_comp_3_T_12 = $signed(w3_mat_comp_3) + $signed(_reg3_mat_comp_3_T_9); // @[calc6x6.scala 154:61]
  wire [37:0] _reg3_mat_comp_9_T_2 = $signed(w3_mat_comp_9) - $signed(w3_mat_comp_15); // @[calc6x6.scala 156:62]
  wire [37:0] _reg3_mat_comp_9_T_5 = $signed(_reg3_mat_comp_9_T_2) + $signed(w3_mat_real_21); // @[calc6x6.scala 156:84]
  wire [37:0] _reg3_mat_comp_9_T_8 = $signed(_reg3_mat_comp_9_T_5) - $signed(w3_mat_real_27); // @[calc6x6.scala 156:106]
  wire [35:0] _GEN_725 = _reg3_mat_comp_9_T_8[37:2]; // @[calc6x6.scala 156:129]
  wire [37:0] _reg3_mat_comp_9_T_9 = {{2{_GEN_725[35]}},_GEN_725}; // @[calc6x6.scala 156:129]
  wire [37:0] _reg3_mat_comp_15_T_5 = $signed(_reg3_mat_comp_3_T_2) - $signed(w3_mat_comp_21); // @[calc6x6.scala 157:84]
  wire [37:0] _reg3_mat_comp_15_T_8 = $signed(_reg3_mat_comp_15_T_5) - $signed(w3_mat_comp_27); // @[calc6x6.scala 157:106]
  wire [35:0] _GEN_726 = _reg3_mat_comp_15_T_8[37:2]; // @[calc6x6.scala 157:129]
  wire [37:0] _reg3_mat_comp_15_T_9 = {{2{_GEN_726[35]}},_GEN_726}; // @[calc6x6.scala 157:129]
  wire [37:0] _reg3_mat_comp_21_T_5 = $signed(_reg3_mat_comp_9_T_2) - $signed(w3_mat_real_21); // @[calc6x6.scala 158:85]
  wire [37:0] _reg3_mat_comp_21_T_8 = $signed(_reg3_mat_comp_21_T_5) + $signed(w3_mat_real_27); // @[calc6x6.scala 158:107]
  wire [35:0] _GEN_727 = _reg3_mat_comp_21_T_8[37:2]; // @[calc6x6.scala 158:130]
  wire [37:0] _reg3_mat_comp_21_T_9 = {{2{_GEN_727[35]}},_GEN_727}; // @[calc6x6.scala 158:130]
  wire [37:0] _reg3_mat_comp_21_T_12 = $signed(_reg3_mat_comp_21_T_9) + $signed(w3_mat_comp_33); // @[calc6x6.scala 158:136]
  wire [37:0] _reg3_mat_real_4_T_2 = $signed(w3_mat_real_10) + $signed(w3_mat_real_16); // @[calc6x6.scala 148:85]
  wire [37:0] _reg3_mat_real_4_T_5 = $signed(_reg3_mat_real_4_T_2) + $signed(w3_mat_real_22); // @[calc6x6.scala 149:62]
  wire [37:0] _reg3_mat_real_4_T_8 = $signed(_reg3_mat_real_4_T_5) + $signed(w3_mat_real_28); // @[calc6x6.scala 149:84]
  wire [35:0] _GEN_728 = _reg3_mat_real_4_T_8[37:2]; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_4_T_9 = {{2{_GEN_728[35]}},_GEN_728}; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_4_T_12 = $signed(w3_mat_real_4) + $signed(_reg3_mat_real_4_T_9); // @[calc6x6.scala 148:61]
  wire [37:0] _reg3_mat_real_10_T_2 = $signed(w3_mat_real_10) - $signed(w3_mat_real_16); // @[calc6x6.scala 150:62]
  wire [37:0] _reg3_mat_real_10_T_5 = $signed(_reg3_mat_real_10_T_2) - $signed(w3_mat_comp_22); // @[calc6x6.scala 150:84]
  wire [37:0] _reg3_mat_real_10_T_8 = $signed(_reg3_mat_real_10_T_5) + $signed(w3_mat_comp_28); // @[calc6x6.scala 150:106]
  wire [35:0] _GEN_729 = _reg3_mat_real_10_T_8[37:2]; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_10_T_9 = {{2{_GEN_729[35]}},_GEN_729}; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_16_T_5 = $signed(_reg3_mat_real_4_T_2) - $signed(w3_mat_real_22); // @[calc6x6.scala 151:84]
  wire [37:0] _reg3_mat_real_16_T_8 = $signed(_reg3_mat_real_16_T_5) - $signed(w3_mat_real_28); // @[calc6x6.scala 151:106]
  wire [35:0] _GEN_730 = _reg3_mat_real_16_T_8[37:2]; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_16_T_9 = {{2{_GEN_730[35]}},_GEN_730}; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_22_T_5 = $signed(_reg3_mat_real_10_T_2) + $signed(w3_mat_comp_22); // @[calc6x6.scala 152:85]
  wire [37:0] _reg3_mat_real_22_T_8 = $signed(_reg3_mat_real_22_T_5) - $signed(w3_mat_comp_28); // @[calc6x6.scala 152:107]
  wire [35:0] _GEN_731 = _reg3_mat_real_22_T_8[37:2]; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_22_T_9 = {{2{_GEN_731[35]}},_GEN_731}; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_22_T_12 = $signed(_reg3_mat_real_22_T_9) + $signed(w3_mat_real_34); // @[calc6x6.scala 152:136]
  wire [37:0] _reg3_mat_comp_4_T_2 = $signed(w3_mat_comp_10) + $signed(w3_mat_comp_16); // @[calc6x6.scala 154:85]
  wire [37:0] _reg3_mat_comp_4_T_5 = $signed(_reg3_mat_comp_4_T_2) + $signed(w3_mat_comp_22); // @[calc6x6.scala 155:62]
  wire [37:0] _reg3_mat_comp_4_T_8 = $signed(_reg3_mat_comp_4_T_5) + $signed(w3_mat_comp_28); // @[calc6x6.scala 155:84]
  wire [35:0] _GEN_732 = _reg3_mat_comp_4_T_8[37:2]; // @[calc6x6.scala 155:107]
  wire [37:0] _reg3_mat_comp_4_T_9 = {{2{_GEN_732[35]}},_GEN_732}; // @[calc6x6.scala 155:107]
  wire [37:0] _reg3_mat_comp_4_T_12 = $signed(w3_mat_comp_4) + $signed(_reg3_mat_comp_4_T_9); // @[calc6x6.scala 154:61]
  wire [37:0] _reg3_mat_comp_10_T_2 = $signed(w3_mat_comp_10) - $signed(w3_mat_comp_16); // @[calc6x6.scala 156:62]
  wire [37:0] _reg3_mat_comp_10_T_5 = $signed(_reg3_mat_comp_10_T_2) + $signed(w3_mat_real_22); // @[calc6x6.scala 156:84]
  wire [37:0] _reg3_mat_comp_10_T_8 = $signed(_reg3_mat_comp_10_T_5) - $signed(w3_mat_real_28); // @[calc6x6.scala 156:106]
  wire [35:0] _GEN_733 = _reg3_mat_comp_10_T_8[37:2]; // @[calc6x6.scala 156:129]
  wire [37:0] _reg3_mat_comp_10_T_9 = {{2{_GEN_733[35]}},_GEN_733}; // @[calc6x6.scala 156:129]
  wire [37:0] _reg3_mat_comp_16_T_5 = $signed(_reg3_mat_comp_4_T_2) - $signed(w3_mat_comp_22); // @[calc6x6.scala 157:84]
  wire [37:0] _reg3_mat_comp_16_T_8 = $signed(_reg3_mat_comp_16_T_5) - $signed(w3_mat_comp_28); // @[calc6x6.scala 157:106]
  wire [35:0] _GEN_734 = _reg3_mat_comp_16_T_8[37:2]; // @[calc6x6.scala 157:129]
  wire [37:0] _reg3_mat_comp_16_T_9 = {{2{_GEN_734[35]}},_GEN_734}; // @[calc6x6.scala 157:129]
  wire [37:0] _reg3_mat_comp_22_T_5 = $signed(_reg3_mat_comp_10_T_2) - $signed(w3_mat_real_22); // @[calc6x6.scala 158:85]
  wire [37:0] _reg3_mat_comp_22_T_8 = $signed(_reg3_mat_comp_22_T_5) + $signed(w3_mat_real_28); // @[calc6x6.scala 158:107]
  wire [35:0] _GEN_735 = _reg3_mat_comp_22_T_8[37:2]; // @[calc6x6.scala 158:130]
  wire [37:0] _reg3_mat_comp_22_T_9 = {{2{_GEN_735[35]}},_GEN_735}; // @[calc6x6.scala 158:130]
  wire [37:0] _reg3_mat_comp_22_T_12 = $signed(_reg3_mat_comp_22_T_9) + $signed(w3_mat_comp_34); // @[calc6x6.scala 158:136]
  wire [37:0] _reg3_mat_real_5_T_2 = $signed(w3_mat_real_11) + $signed(w3_mat_real_17); // @[calc6x6.scala 148:85]
  wire [37:0] _reg3_mat_real_5_T_5 = $signed(_reg3_mat_real_5_T_2) + $signed(w3_mat_real_23); // @[calc6x6.scala 149:62]
  wire [37:0] _reg3_mat_real_5_T_8 = $signed(_reg3_mat_real_5_T_5) + $signed(w3_mat_real_29); // @[calc6x6.scala 149:84]
  wire [35:0] _GEN_736 = _reg3_mat_real_5_T_8[37:2]; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_5_T_9 = {{2{_GEN_736[35]}},_GEN_736}; // @[calc6x6.scala 149:107]
  wire [37:0] _reg3_mat_real_5_T_12 = $signed(w3_mat_real_5) + $signed(_reg3_mat_real_5_T_9); // @[calc6x6.scala 148:61]
  wire [37:0] _reg3_mat_real_11_T_2 = $signed(w3_mat_real_11) - $signed(w3_mat_real_17); // @[calc6x6.scala 150:62]
  wire [37:0] _reg3_mat_real_11_T_5 = $signed(_reg3_mat_real_11_T_2) - $signed(w3_mat_comp_23); // @[calc6x6.scala 150:84]
  wire [37:0] _reg3_mat_real_11_T_8 = $signed(_reg3_mat_real_11_T_5) + $signed(w3_mat_comp_29); // @[calc6x6.scala 150:106]
  wire [35:0] _GEN_737 = _reg3_mat_real_11_T_8[37:2]; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_11_T_9 = {{2{_GEN_737[35]}},_GEN_737}; // @[calc6x6.scala 150:129]
  wire [37:0] _reg3_mat_real_17_T_5 = $signed(_reg3_mat_real_5_T_2) - $signed(w3_mat_real_23); // @[calc6x6.scala 151:84]
  wire [37:0] _reg3_mat_real_17_T_8 = $signed(_reg3_mat_real_17_T_5) - $signed(w3_mat_real_29); // @[calc6x6.scala 151:106]
  wire [35:0] _GEN_738 = _reg3_mat_real_17_T_8[37:2]; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_17_T_9 = {{2{_GEN_738[35]}},_GEN_738}; // @[calc6x6.scala 151:129]
  wire [37:0] _reg3_mat_real_23_T_5 = $signed(_reg3_mat_real_11_T_2) + $signed(w3_mat_comp_23); // @[calc6x6.scala 152:85]
  wire [37:0] _reg3_mat_real_23_T_8 = $signed(_reg3_mat_real_23_T_5) - $signed(w3_mat_comp_29); // @[calc6x6.scala 152:107]
  wire [35:0] _GEN_739 = _reg3_mat_real_23_T_8[37:2]; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_23_T_9 = {{2{_GEN_739[35]}},_GEN_739}; // @[calc6x6.scala 152:130]
  wire [37:0] _reg3_mat_real_23_T_12 = $signed(_reg3_mat_real_23_T_9) + $signed(w3_mat_real_35); // @[calc6x6.scala 152:136]
  wire  _T_2 = 2'h0 == io_flag; // @[Conditional.scala 37:30]
  wire  _T_5 = 2'h1 == io_flag; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h2 == io_flag; // @[Conditional.scala 37:30]
  wire [37:0] _io_output_mat_0_T_2 = $signed(reg3_mat_real_1) + $signed(reg3_mat_real_2); // @[calc6x6.scala 164:85]
  wire [37:0] _io_output_mat_0_T_5 = $signed(_io_output_mat_0_T_2) + $signed(reg3_mat_real_3); // @[calc6x6.scala 165:62]
  wire [37:0] _io_output_mat_0_T_8 = $signed(_io_output_mat_0_T_5) + $signed(reg3_mat_real_4); // @[calc6x6.scala 165:84]
  wire [35:0] _GEN_744 = _io_output_mat_0_T_8[37:2]; // @[calc6x6.scala 165:107]
  wire [37:0] _io_output_mat_0_T_9 = {{2{_GEN_744[35]}},_GEN_744}; // @[calc6x6.scala 165:107]
  wire [37:0] _io_output_mat_0_T_12 = $signed(reg3_mat_real_0) + $signed(_io_output_mat_0_T_9); // @[calc6x6.scala 164:61]
  wire [37:0] _io_output_mat_1_T_2 = $signed(reg3_mat_real_1) - $signed(reg3_mat_real_2); // @[calc6x6.scala 166:63]
  wire [37:0] _io_output_mat_1_T_5 = $signed(_io_output_mat_1_T_2) - $signed(reg3_mat_comp_3); // @[calc6x6.scala 166:85]
  wire [37:0] _io_output_mat_1_T_8 = $signed(_io_output_mat_1_T_5) + $signed(reg3_mat_comp_4); // @[calc6x6.scala 166:107]
  wire [35:0] _GEN_745 = _io_output_mat_1_T_8[37:2]; // @[calc6x6.scala 166:130]
  wire [37:0] _io_output_mat_1_T_9 = {{2{_GEN_745[35]}},_GEN_745}; // @[calc6x6.scala 166:130]
  wire [37:0] _io_output_mat_2_T_5 = $signed(_io_output_mat_0_T_2) - $signed(reg3_mat_real_3); // @[calc6x6.scala 167:85]
  wire [37:0] _io_output_mat_2_T_8 = $signed(_io_output_mat_2_T_5) - $signed(reg3_mat_real_4); // @[calc6x6.scala 167:107]
  wire [35:0] _GEN_746 = _io_output_mat_2_T_8[37:2]; // @[calc6x6.scala 167:130]
  wire [37:0] _io_output_mat_2_T_9 = {{2{_GEN_746[35]}},_GEN_746}; // @[calc6x6.scala 167:130]
  wire [37:0] _io_output_mat_3_T_5 = $signed(_io_output_mat_1_T_2) + $signed(reg3_mat_comp_3); // @[calc6x6.scala 168:85]
  wire [37:0] _io_output_mat_3_T_8 = $signed(_io_output_mat_3_T_5) - $signed(reg3_mat_comp_4); // @[calc6x6.scala 168:107]
  wire [35:0] _GEN_747 = _io_output_mat_3_T_8[37:2]; // @[calc6x6.scala 168:130]
  wire [37:0] _io_output_mat_3_T_9 = {{2{_GEN_747[35]}},_GEN_747}; // @[calc6x6.scala 168:130]
  wire [37:0] _io_output_mat_3_T_12 = $signed(_io_output_mat_3_T_9) + $signed(reg3_mat_real_5); // @[calc6x6.scala 168:136]
  wire [37:0] _io_output_mat_4_T_2 = $signed(reg3_mat_real_7) + $signed(reg3_mat_real_8); // @[calc6x6.scala 164:85]
  wire [37:0] _io_output_mat_4_T_5 = $signed(_io_output_mat_4_T_2) + $signed(reg3_mat_real_9); // @[calc6x6.scala 165:62]
  wire [37:0] _io_output_mat_4_T_8 = $signed(_io_output_mat_4_T_5) + $signed(reg3_mat_real_10); // @[calc6x6.scala 165:84]
  wire [35:0] _GEN_748 = _io_output_mat_4_T_8[37:2]; // @[calc6x6.scala 165:107]
  wire [37:0] _io_output_mat_4_T_9 = {{2{_GEN_748[35]}},_GEN_748}; // @[calc6x6.scala 165:107]
  wire [37:0] _io_output_mat_4_T_12 = $signed(reg3_mat_real_6) + $signed(_io_output_mat_4_T_9); // @[calc6x6.scala 164:61]
  wire [37:0] _io_output_mat_5_T_2 = $signed(reg3_mat_real_7) - $signed(reg3_mat_real_8); // @[calc6x6.scala 166:63]
  wire [37:0] _io_output_mat_5_T_5 = $signed(_io_output_mat_5_T_2) - $signed(reg3_mat_comp_9); // @[calc6x6.scala 166:85]
  wire [37:0] _io_output_mat_5_T_8 = $signed(_io_output_mat_5_T_5) + $signed(reg3_mat_comp_10); // @[calc6x6.scala 166:107]
  wire [35:0] _GEN_749 = _io_output_mat_5_T_8[37:2]; // @[calc6x6.scala 166:130]
  wire [37:0] _io_output_mat_5_T_9 = {{2{_GEN_749[35]}},_GEN_749}; // @[calc6x6.scala 166:130]
  wire [37:0] _io_output_mat_6_T_5 = $signed(_io_output_mat_4_T_2) - $signed(reg3_mat_real_9); // @[calc6x6.scala 167:85]
  wire [37:0] _io_output_mat_6_T_8 = $signed(_io_output_mat_6_T_5) - $signed(reg3_mat_real_10); // @[calc6x6.scala 167:107]
  wire [35:0] _GEN_750 = _io_output_mat_6_T_8[37:2]; // @[calc6x6.scala 167:130]
  wire [37:0] _io_output_mat_6_T_9 = {{2{_GEN_750[35]}},_GEN_750}; // @[calc6x6.scala 167:130]
  wire [37:0] _io_output_mat_7_T_5 = $signed(_io_output_mat_5_T_2) + $signed(reg3_mat_comp_9); // @[calc6x6.scala 168:85]
  wire [37:0] _io_output_mat_7_T_8 = $signed(_io_output_mat_7_T_5) - $signed(reg3_mat_comp_10); // @[calc6x6.scala 168:107]
  wire [35:0] _GEN_751 = _io_output_mat_7_T_8[37:2]; // @[calc6x6.scala 168:130]
  wire [37:0] _io_output_mat_7_T_9 = {{2{_GEN_751[35]}},_GEN_751}; // @[calc6x6.scala 168:130]
  wire [37:0] _io_output_mat_7_T_12 = $signed(_io_output_mat_7_T_9) + $signed(reg3_mat_real_11); // @[calc6x6.scala 168:136]
  wire [37:0] _io_output_mat_8_T_2 = $signed(reg3_mat_real_13) + $signed(reg3_mat_real_14); // @[calc6x6.scala 164:85]
  wire [37:0] _io_output_mat_8_T_5 = $signed(_io_output_mat_8_T_2) + $signed(reg3_mat_real_15); // @[calc6x6.scala 165:62]
  wire [37:0] _io_output_mat_8_T_8 = $signed(_io_output_mat_8_T_5) + $signed(reg3_mat_real_16); // @[calc6x6.scala 165:84]
  wire [35:0] _GEN_752 = _io_output_mat_8_T_8[37:2]; // @[calc6x6.scala 165:107]
  wire [37:0] _io_output_mat_8_T_9 = {{2{_GEN_752[35]}},_GEN_752}; // @[calc6x6.scala 165:107]
  wire [37:0] _io_output_mat_8_T_12 = $signed(reg3_mat_real_12) + $signed(_io_output_mat_8_T_9); // @[calc6x6.scala 164:61]
  wire [37:0] _io_output_mat_9_T_2 = $signed(reg3_mat_real_13) - $signed(reg3_mat_real_14); // @[calc6x6.scala 166:63]
  wire [37:0] _io_output_mat_9_T_5 = $signed(_io_output_mat_9_T_2) - $signed(reg3_mat_comp_15); // @[calc6x6.scala 166:85]
  wire [37:0] _io_output_mat_9_T_8 = $signed(_io_output_mat_9_T_5) + $signed(reg3_mat_comp_16); // @[calc6x6.scala 166:107]
  wire [35:0] _GEN_753 = _io_output_mat_9_T_8[37:2]; // @[calc6x6.scala 166:130]
  wire [37:0] _io_output_mat_9_T_9 = {{2{_GEN_753[35]}},_GEN_753}; // @[calc6x6.scala 166:130]
  wire [37:0] _io_output_mat_10_T_5 = $signed(_io_output_mat_8_T_2) - $signed(reg3_mat_real_15); // @[calc6x6.scala 167:85]
  wire [37:0] _io_output_mat_10_T_8 = $signed(_io_output_mat_10_T_5) - $signed(reg3_mat_real_16); // @[calc6x6.scala 167:107]
  wire [35:0] _GEN_754 = _io_output_mat_10_T_8[37:2]; // @[calc6x6.scala 167:130]
  wire [37:0] _io_output_mat_10_T_9 = {{2{_GEN_754[35]}},_GEN_754}; // @[calc6x6.scala 167:130]
  wire [37:0] _io_output_mat_11_T_5 = $signed(_io_output_mat_9_T_2) + $signed(reg3_mat_comp_15); // @[calc6x6.scala 168:85]
  wire [37:0] _io_output_mat_11_T_8 = $signed(_io_output_mat_11_T_5) - $signed(reg3_mat_comp_16); // @[calc6x6.scala 168:107]
  wire [35:0] _GEN_755 = _io_output_mat_11_T_8[37:2]; // @[calc6x6.scala 168:130]
  wire [37:0] _io_output_mat_11_T_9 = {{2{_GEN_755[35]}},_GEN_755}; // @[calc6x6.scala 168:130]
  wire [37:0] _io_output_mat_11_T_12 = $signed(_io_output_mat_11_T_9) + $signed(reg3_mat_real_17); // @[calc6x6.scala 168:136]
  wire [37:0] _io_output_mat_12_T_2 = $signed(reg3_mat_real_19) + $signed(reg3_mat_real_20); // @[calc6x6.scala 164:85]
  wire [37:0] _io_output_mat_12_T_5 = $signed(_io_output_mat_12_T_2) + $signed(reg3_mat_real_21); // @[calc6x6.scala 165:62]
  wire [37:0] _io_output_mat_12_T_8 = $signed(_io_output_mat_12_T_5) + $signed(reg3_mat_real_22); // @[calc6x6.scala 165:84]
  wire [35:0] _GEN_756 = _io_output_mat_12_T_8[37:2]; // @[calc6x6.scala 165:107]
  wire [37:0] _io_output_mat_12_T_9 = {{2{_GEN_756[35]}},_GEN_756}; // @[calc6x6.scala 165:107]
  wire [37:0] _io_output_mat_12_T_12 = $signed(reg3_mat_real_18) + $signed(_io_output_mat_12_T_9); // @[calc6x6.scala 164:61]
  wire [37:0] _io_output_mat_13_T_2 = $signed(reg3_mat_real_19) - $signed(reg3_mat_real_20); // @[calc6x6.scala 166:63]
  wire [37:0] _io_output_mat_13_T_5 = $signed(_io_output_mat_13_T_2) - $signed(reg3_mat_comp_21); // @[calc6x6.scala 166:85]
  wire [37:0] _io_output_mat_13_T_8 = $signed(_io_output_mat_13_T_5) + $signed(reg3_mat_comp_22); // @[calc6x6.scala 166:107]
  wire [35:0] _GEN_757 = _io_output_mat_13_T_8[37:2]; // @[calc6x6.scala 166:130]
  wire [37:0] _io_output_mat_13_T_9 = {{2{_GEN_757[35]}},_GEN_757}; // @[calc6x6.scala 166:130]
  wire [37:0] _io_output_mat_14_T_5 = $signed(_io_output_mat_12_T_2) - $signed(reg3_mat_real_21); // @[calc6x6.scala 167:85]
  wire [37:0] _io_output_mat_14_T_8 = $signed(_io_output_mat_14_T_5) - $signed(reg3_mat_real_22); // @[calc6x6.scala 167:107]
  wire [35:0] _GEN_758 = _io_output_mat_14_T_8[37:2]; // @[calc6x6.scala 167:130]
  wire [37:0] _io_output_mat_14_T_9 = {{2{_GEN_758[35]}},_GEN_758}; // @[calc6x6.scala 167:130]
  wire [37:0] _io_output_mat_15_T_5 = $signed(_io_output_mat_13_T_2) + $signed(reg3_mat_comp_21); // @[calc6x6.scala 168:85]
  wire [37:0] _io_output_mat_15_T_8 = $signed(_io_output_mat_15_T_5) - $signed(reg3_mat_comp_22); // @[calc6x6.scala 168:107]
  wire [35:0] _GEN_759 = _io_output_mat_15_T_8[37:2]; // @[calc6x6.scala 168:130]
  wire [37:0] _io_output_mat_15_T_9 = {{2{_GEN_759[35]}},_GEN_759}; // @[calc6x6.scala 168:130]
  wire [37:0] _io_output_mat_15_T_12 = $signed(_io_output_mat_15_T_9) + $signed(reg3_mat_real_23); // @[calc6x6.scala 168:136]
  wire [19:0] _comp1_0_in_b_T_3 = $signed(reg2_mat_real_3) + $signed(reg2_mat_comp_6); // @[calc6x6.scala 261:65]
  wire [42:0] comp2_0_result = Core_26_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_0_result = Core_36_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_3_T_2 = $signed(comp2_0_result) - $signed(comp3_0_result); // @[calc6x6.scala 264:65]
  wire [42:0] comp1_0_result = Core_16_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_3_T_2 = $signed(comp1_0_result) - $signed(comp2_0_result); // @[calc6x6.scala 265:65]
  wire [42:0] _w3_mat_comp_3_T_5 = $signed(_w3_mat_comp_3_T_2) - $signed(comp3_0_result); // @[calc6x6.scala 265:81]
  wire [42:0] _w3_mat_comp_4_T_2 = 43'sh0 - $signed(comp1_0_result); // @[calc6x6.scala 272:50]
  wire [42:0] _w3_mat_comp_4_T_5 = $signed(_w3_mat_comp_4_T_2) + $signed(comp2_0_result); // @[calc6x6.scala 272:71]
  wire [42:0] _w3_mat_comp_4_T_8 = $signed(_w3_mat_comp_4_T_5) + $signed(comp3_0_result); // @[calc6x6.scala 272:92]
  wire [19:0] _comp1_1_in_b_T_3 = $signed(reg2_mat_real_9) + $signed(reg2_mat_comp_7); // @[calc6x6.scala 261:65]
  wire [42:0] comp2_1_result = Core_27_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_1_result = Core_37_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_9_T_2 = $signed(comp2_1_result) - $signed(comp3_1_result); // @[calc6x6.scala 264:65]
  wire [42:0] comp1_1_result = Core_17_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_9_T_2 = $signed(comp1_1_result) - $signed(comp2_1_result); // @[calc6x6.scala 265:65]
  wire [42:0] _w3_mat_comp_9_T_5 = $signed(_w3_mat_comp_9_T_2) - $signed(comp3_1_result); // @[calc6x6.scala 265:81]
  wire [42:0] _w3_mat_comp_10_T_2 = 43'sh0 - $signed(comp1_1_result); // @[calc6x6.scala 272:50]
  wire [42:0] _w3_mat_comp_10_T_5 = $signed(_w3_mat_comp_10_T_2) + $signed(comp2_1_result); // @[calc6x6.scala 272:71]
  wire [42:0] _w3_mat_comp_10_T_8 = $signed(_w3_mat_comp_10_T_5) + $signed(comp3_1_result); // @[calc6x6.scala 272:92]
  wire [19:0] _comp1_2_in_b_T_3 = $signed(reg2_mat_real_15) + $signed(reg2_mat_comp_8); // @[calc6x6.scala 261:65]
  wire [42:0] comp2_2_result = Core_28_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_2_result = Core_38_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_15_T_2 = $signed(comp2_2_result) - $signed(comp3_2_result); // @[calc6x6.scala 264:65]
  wire [42:0] comp1_2_result = Core_18_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_15_T_2 = $signed(comp1_2_result) - $signed(comp2_2_result); // @[calc6x6.scala 265:65]
  wire [42:0] _w3_mat_comp_15_T_5 = $signed(_w3_mat_comp_15_T_2) - $signed(comp3_2_result); // @[calc6x6.scala 265:81]
  wire [42:0] _w3_mat_comp_16_T_2 = 43'sh0 - $signed(comp1_2_result); // @[calc6x6.scala 272:50]
  wire [42:0] _w3_mat_comp_16_T_5 = $signed(_w3_mat_comp_16_T_2) + $signed(comp2_2_result); // @[calc6x6.scala 272:71]
  wire [42:0] _w3_mat_comp_16_T_8 = $signed(_w3_mat_comp_16_T_5) + $signed(comp3_2_result); // @[calc6x6.scala 272:92]
  wire [19:0] _comp1_3_in_b_T_3 = $signed(reg2_mat_real_18) + $signed(reg2_mat_comp_0); // @[calc6x6.scala 238:65]
  wire [42:0] comp2_3_result = Core_29_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_3_result = Core_39_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_18_T_2 = $signed(comp2_3_result) - $signed(comp3_3_result); // @[calc6x6.scala 241:65]
  wire [42:0] comp1_3_result = Core_19_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_18_T_2 = $signed(comp1_3_result) - $signed(comp2_3_result); // @[calc6x6.scala 242:65]
  wire [42:0] _w3_mat_comp_18_T_5 = $signed(_w3_mat_comp_18_T_2) - $signed(comp3_3_result); // @[calc6x6.scala 242:81]
  wire [19:0] _comp1_4_in_b_T_3 = $signed(reg2_mat_real_19) + $signed(reg2_mat_comp_1); // @[calc6x6.scala 238:65]
  wire [42:0] comp2_4_result = Core_30_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_4_result = Core_40_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_19_T_2 = $signed(comp2_4_result) - $signed(comp3_4_result); // @[calc6x6.scala 241:65]
  wire [42:0] comp1_4_result = Core_20_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_19_T_2 = $signed(comp1_4_result) - $signed(comp2_4_result); // @[calc6x6.scala 242:65]
  wire [42:0] _w3_mat_comp_19_T_5 = $signed(_w3_mat_comp_19_T_2) - $signed(comp3_4_result); // @[calc6x6.scala 242:81]
  wire [19:0] _comp1_5_in_b_T_3 = $signed(reg2_mat_real_20) + $signed(reg2_mat_comp_2); // @[calc6x6.scala 238:65]
  wire [42:0] comp2_5_result = Core_31_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_5_result = Core_41_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_20_T_2 = $signed(comp2_5_result) - $signed(comp3_5_result); // @[calc6x6.scala 241:65]
  wire [42:0] comp1_5_result = Core_21_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_20_T_2 = $signed(comp1_5_result) - $signed(comp2_5_result); // @[calc6x6.scala 242:65]
  wire [42:0] _w3_mat_comp_20_T_5 = $signed(_w3_mat_comp_20_T_2) - $signed(comp3_5_result); // @[calc6x6.scala 242:81]
  wire [19:0] _comp1_6_in_b_T_3 = $signed(reg2_mat_real_21) + $signed(reg2_mat_comp_3); // @[calc6x6.scala 238:65]
  wire [42:0] comp2_6_result = Core_32_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_6_result = Core_42_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_21_T_2 = $signed(comp2_6_result) - $signed(comp3_6_result); // @[calc6x6.scala 241:65]
  wire [42:0] comp1_6_result = Core_22_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_21_T_2 = $signed(comp1_6_result) - $signed(comp2_6_result); // @[calc6x6.scala 242:65]
  wire [42:0] _w3_mat_comp_21_T_5 = $signed(_w3_mat_comp_21_T_2) - $signed(comp3_6_result); // @[calc6x6.scala 242:81]
  wire [19:0] _comp1_7_in_b_T_3 = $signed(reg2_mat_real_22) + $signed(reg2_mat_comp_4); // @[calc6x6.scala 238:65]
  wire [42:0] comp2_7_result = Core_33_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_7_result = Core_43_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_22_T_2 = $signed(comp2_7_result) - $signed(comp3_7_result); // @[calc6x6.scala 241:65]
  wire [42:0] comp1_7_result = Core_23_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_22_T_2 = $signed(comp1_7_result) - $signed(comp2_7_result); // @[calc6x6.scala 242:65]
  wire [42:0] _w3_mat_comp_22_T_5 = $signed(_w3_mat_comp_22_T_2) - $signed(comp3_7_result); // @[calc6x6.scala 242:81]
  wire [19:0] _comp1_8_in_b_T_3 = $signed(reg2_mat_real_23) + $signed(reg2_mat_comp_5); // @[calc6x6.scala 238:65]
  wire [42:0] comp2_8_result = Core_34_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_8_result = Core_44_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_23_T_2 = $signed(comp2_8_result) - $signed(comp3_8_result); // @[calc6x6.scala 241:65]
  wire [42:0] comp1_8_result = Core_24_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_23_T_2 = $signed(comp1_8_result) - $signed(comp2_8_result); // @[calc6x6.scala 242:65]
  wire [42:0] _w3_mat_comp_23_T_5 = $signed(_w3_mat_comp_23_T_2) - $signed(comp3_8_result); // @[calc6x6.scala 242:81]
  wire [42:0] _w3_mat_comp_24_T_2 = 43'sh0 - $signed(comp1_3_result); // @[calc6x6.scala 250:50]
  wire [42:0] _w3_mat_comp_24_T_5 = $signed(_w3_mat_comp_24_T_2) + $signed(comp2_3_result); // @[calc6x6.scala 250:71]
  wire [42:0] _w3_mat_comp_24_T_8 = $signed(_w3_mat_comp_24_T_5) + $signed(comp3_3_result); // @[calc6x6.scala 250:92]
  wire [42:0] _w3_mat_comp_25_T_2 = 43'sh0 - $signed(comp1_4_result); // @[calc6x6.scala 250:50]
  wire [42:0] _w3_mat_comp_25_T_5 = $signed(_w3_mat_comp_25_T_2) + $signed(comp2_4_result); // @[calc6x6.scala 250:71]
  wire [42:0] _w3_mat_comp_25_T_8 = $signed(_w3_mat_comp_25_T_5) + $signed(comp3_4_result); // @[calc6x6.scala 250:92]
  wire [42:0] _w3_mat_comp_26_T_2 = 43'sh0 - $signed(comp1_5_result); // @[calc6x6.scala 250:50]
  wire [42:0] _w3_mat_comp_26_T_5 = $signed(_w3_mat_comp_26_T_2) + $signed(comp2_5_result); // @[calc6x6.scala 250:71]
  wire [42:0] _w3_mat_comp_26_T_8 = $signed(_w3_mat_comp_26_T_5) + $signed(comp3_5_result); // @[calc6x6.scala 250:92]
  wire [42:0] _w3_mat_comp_27_T_2 = 43'sh0 - $signed(comp1_7_result); // @[calc6x6.scala 250:50]
  wire [42:0] _w3_mat_comp_27_T_5 = $signed(_w3_mat_comp_27_T_2) + $signed(comp2_7_result); // @[calc6x6.scala 250:71]
  wire [42:0] _w3_mat_comp_27_T_8 = $signed(_w3_mat_comp_27_T_5) + $signed(comp3_7_result); // @[calc6x6.scala 250:92]
  wire [42:0] _w3_mat_comp_28_T_2 = 43'sh0 - $signed(comp1_6_result); // @[calc6x6.scala 250:50]
  wire [42:0] _w3_mat_comp_28_T_5 = $signed(_w3_mat_comp_28_T_2) + $signed(comp2_6_result); // @[calc6x6.scala 250:71]
  wire [42:0] _w3_mat_comp_28_T_8 = $signed(_w3_mat_comp_28_T_5) + $signed(comp3_6_result); // @[calc6x6.scala 250:92]
  wire [42:0] _w3_mat_comp_29_T_2 = 43'sh0 - $signed(comp1_8_result); // @[calc6x6.scala 250:50]
  wire [42:0] _w3_mat_comp_29_T_5 = $signed(_w3_mat_comp_29_T_2) + $signed(comp2_8_result); // @[calc6x6.scala 250:71]
  wire [42:0] _w3_mat_comp_29_T_8 = $signed(_w3_mat_comp_29_T_5) + $signed(comp3_8_result); // @[calc6x6.scala 250:92]
  wire [19:0] _comp1_9_in_b_T_3 = $signed(reg2_mat_real_33) + $signed(reg2_mat_comp_9); // @[calc6x6.scala 261:65]
  wire [42:0] comp2_9_result = Core_35_io_result; // @[calc6x6.scala 72:24 calc6x6.scala 72:24]
  wire [42:0] comp3_9_result = Core_45_io_result; // @[calc6x6.scala 73:24 calc6x6.scala 73:24]
  wire [42:0] _w3_mat_real_33_T_2 = $signed(comp2_9_result) - $signed(comp3_9_result); // @[calc6x6.scala 264:65]
  wire [42:0] comp1_9_result = Core_25_io_result; // @[calc6x6.scala 71:24 calc6x6.scala 71:24]
  wire [42:0] _w3_mat_comp_33_T_2 = $signed(comp1_9_result) - $signed(comp2_9_result); // @[calc6x6.scala 265:65]
  wire [42:0] _w3_mat_comp_33_T_5 = $signed(_w3_mat_comp_33_T_2) - $signed(comp3_9_result); // @[calc6x6.scala 265:81]
  wire [42:0] _w3_mat_comp_34_T_2 = 43'sh0 - $signed(comp1_9_result); // @[calc6x6.scala 272:50]
  wire [42:0] _w3_mat_comp_34_T_5 = $signed(_w3_mat_comp_34_T_2) + $signed(comp2_9_result); // @[calc6x6.scala 272:71]
  wire [42:0] _w3_mat_comp_34_T_8 = $signed(_w3_mat_comp_34_T_5) + $signed(comp3_9_result); // @[calc6x6.scala 272:92]
  wire [37:0] _GEN_0 = _T_8 ? $signed(_io_output_mat_0_T_12) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 164:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_1 = _T_8 ? $signed(_io_output_mat_1_T_9) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 166:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_2 = _T_8 ? $signed(_io_output_mat_2_T_9) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 167:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_3 = _T_8 ? $signed(_io_output_mat_3_T_12) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 168:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_4 = _T_8 ? $signed(_io_output_mat_4_T_12) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 164:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_5 = _T_8 ? $signed(_io_output_mat_5_T_9) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 166:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_6 = _T_8 ? $signed(_io_output_mat_6_T_9) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 167:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_7 = _T_8 ? $signed(_io_output_mat_7_T_12) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 168:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_8 = _T_8 ? $signed(_io_output_mat_8_T_12) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 164:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_9 = _T_8 ? $signed(_io_output_mat_9_T_9) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 166:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_10 = _T_8 ? $signed(_io_output_mat_10_T_9) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 167:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_11 = _T_8 ? $signed(_io_output_mat_11_T_12) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 168:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_12 = _T_8 ? $signed(_io_output_mat_12_T_12) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 164:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_13 = _T_8 ? $signed(_io_output_mat_13_T_9) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 166:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_14 = _T_8 ? $signed(_io_output_mat_14_T_9) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 167:37 calc6x6.scala 87:15]
  wire [37:0] _GEN_15 = _T_8 ? $signed(_io_output_mat_15_T_12) : $signed(38'sh0); // @[Conditional.scala 39:67 calc6x6.scala 168:37 calc6x6.scala 87:15]
  wire [24:0] _GEN_17 = _T_8 ? $signed({{5{reg2_mat_real_0[19]}},reg2_mat_real_0}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_18 = _T_8 ? $signed(io_weight_real_0) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_0_result = Core_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_19 = _T_8 ? $signed(real_0_result) : $signed({{5{w3_mat_real_0[37]}},w3_mat_real_0}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_21 = _T_8 ? $signed({{5{reg2_mat_real_1[19]}},reg2_mat_real_1}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_22 = _T_8 ? $signed(io_weight_real_1) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_1_result = Core_1_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_23 = _T_8 ? $signed(real_1_result) : $signed({{5{w3_mat_real_1[37]}},w3_mat_real_1}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_25 = _T_8 ? $signed({{5{reg2_mat_real_2[19]}},reg2_mat_real_2}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_26 = _T_8 ? $signed(io_weight_real_2) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_2_result = Core_2_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_27 = _T_8 ? $signed(real_2_result) : $signed({{5{w3_mat_real_2[37]}},w3_mat_real_2}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_31 = _T_8 ? $signed(io_weight_comp1_0) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 257:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_32 = _T_8 ? $signed(io_weight_comp2_0) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 258:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_33 = _T_8 ? $signed(io_weight_comp3_0) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 259:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_34 = _T_8 ? $signed({{5{_comp1_0_in_b_T_3[19]}},_comp1_0_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 261:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_35 = _T_8 ? $signed({{5{reg2_mat_real_3[19]}},reg2_mat_real_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 262:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_36 = _T_8 ? $signed({{5{reg2_mat_comp_6[19]}},reg2_mat_comp_6}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 263:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_37 = _T_8 ? $signed(_w3_mat_real_3_T_2) : $signed({{5{w3_mat_real_3[37]}},w3_mat_real_3}); // @[Conditional.scala 39:67 calc6x6.scala 264:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_38 = _T_8 ? $signed(_w3_mat_comp_3_T_5) : $signed({{5{w3_mat_comp_3[37]}},w3_mat_comp_3}); // @[Conditional.scala 39:67 calc6x6.scala 265:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_39 = _T_8 ? $signed(_w3_mat_real_3_T_2) : $signed({{5{w3_mat_real_4[37]}},w3_mat_real_4}); // @[Conditional.scala 39:67 calc6x6.scala 271:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_40 = _T_8 ? $signed(_w3_mat_comp_4_T_8) : $signed({{5{w3_mat_comp_4[37]}},w3_mat_comp_4}); // @[Conditional.scala 39:67 calc6x6.scala 272:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_42 = _T_8 ? $signed({{5{reg2_mat_real_5[19]}},reg2_mat_real_5}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_43 = _T_8 ? $signed(io_weight_real_3) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_3_result = Core_3_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_44 = _T_8 ? $signed(real_3_result) : $signed({{5{w3_mat_real_5[37]}},w3_mat_real_5}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_46 = _T_8 ? $signed({{5{reg2_mat_real_6[19]}},reg2_mat_real_6}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_47 = _T_8 ? $signed(io_weight_real_4) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_4_result = Core_4_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_48 = _T_8 ? $signed(real_4_result) : $signed({{5{w3_mat_real_6[37]}},w3_mat_real_6}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_50 = _T_8 ? $signed({{5{reg2_mat_real_7[19]}},reg2_mat_real_7}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_51 = _T_8 ? $signed(io_weight_real_5) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_5_result = Core_5_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_52 = _T_8 ? $signed(real_5_result) : $signed({{5{w3_mat_real_7[37]}},w3_mat_real_7}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_54 = _T_8 ? $signed({{5{reg2_mat_real_8[19]}},reg2_mat_real_8}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_55 = _T_8 ? $signed(io_weight_real_6) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_6_result = Core_6_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_56 = _T_8 ? $signed(real_6_result) : $signed({{5{w3_mat_real_8[37]}},w3_mat_real_8}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_60 = _T_8 ? $signed(io_weight_comp1_1) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 257:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_61 = _T_8 ? $signed(io_weight_comp2_1) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 258:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_62 = _T_8 ? $signed(io_weight_comp3_1) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 259:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_63 = _T_8 ? $signed({{5{_comp1_1_in_b_T_3[19]}},_comp1_1_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 261:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_64 = _T_8 ? $signed({{5{reg2_mat_real_9[19]}},reg2_mat_real_9}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 262:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_65 = _T_8 ? $signed({{5{reg2_mat_comp_7[19]}},reg2_mat_comp_7}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 263:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_66 = _T_8 ? $signed(_w3_mat_real_9_T_2) : $signed({{5{w3_mat_real_9[37]}},w3_mat_real_9}); // @[Conditional.scala 39:67 calc6x6.scala 264:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_67 = _T_8 ? $signed(_w3_mat_comp_9_T_5) : $signed({{5{w3_mat_comp_9[37]}},w3_mat_comp_9}); // @[Conditional.scala 39:67 calc6x6.scala 265:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_68 = _T_8 ? $signed(_w3_mat_real_9_T_2) : $signed({{5{w3_mat_real_10[37]}},w3_mat_real_10}); // @[Conditional.scala 39:67 calc6x6.scala 271:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_69 = _T_8 ? $signed(_w3_mat_comp_10_T_8) : $signed({{5{w3_mat_comp_10[37]}},w3_mat_comp_10}); // @[Conditional.scala 39:67 calc6x6.scala 272:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_71 = _T_8 ? $signed({{5{reg2_mat_real_11[19]}},reg2_mat_real_11}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_72 = _T_8 ? $signed(io_weight_real_7) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_7_result = Core_7_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_73 = _T_8 ? $signed(real_7_result) : $signed({{5{w3_mat_real_11[37]}},w3_mat_real_11}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_75 = _T_8 ? $signed({{5{reg2_mat_real_12[19]}},reg2_mat_real_12}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_76 = _T_8 ? $signed(io_weight_real_8) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_8_result = Core_8_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_77 = _T_8 ? $signed(real_8_result) : $signed({{5{w3_mat_real_12[37]}},w3_mat_real_12}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_79 = _T_8 ? $signed({{5{reg2_mat_real_13[19]}},reg2_mat_real_13}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_80 = _T_8 ? $signed(io_weight_real_9) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_9_result = Core_9_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_81 = _T_8 ? $signed(real_9_result) : $signed({{5{w3_mat_real_13[37]}},w3_mat_real_13}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_83 = _T_8 ? $signed({{5{reg2_mat_real_14[19]}},reg2_mat_real_14}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_84 = _T_8 ? $signed(io_weight_real_10) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_10_result = Core_10_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_85 = _T_8 ? $signed(real_10_result) : $signed({{5{w3_mat_real_14[37]}},w3_mat_real_14}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_89 = _T_8 ? $signed(io_weight_comp1_2) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 257:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_90 = _T_8 ? $signed(io_weight_comp2_2) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 258:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_91 = _T_8 ? $signed(io_weight_comp3_2) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 259:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_92 = _T_8 ? $signed({{5{_comp1_2_in_b_T_3[19]}},_comp1_2_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 261:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_93 = _T_8 ? $signed({{5{reg2_mat_real_15[19]}},reg2_mat_real_15}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 262:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_94 = _T_8 ? $signed({{5{reg2_mat_comp_8[19]}},reg2_mat_comp_8}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 263:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_95 = _T_8 ? $signed(_w3_mat_real_15_T_2) : $signed({{5{w3_mat_real_15[37]}},w3_mat_real_15}); // @[Conditional.scala 39:67 calc6x6.scala 264:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_96 = _T_8 ? $signed(_w3_mat_comp_15_T_5) : $signed({{5{w3_mat_comp_15[37]}},w3_mat_comp_15}); // @[Conditional.scala 39:67 calc6x6.scala 265:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_97 = _T_8 ? $signed(_w3_mat_real_15_T_2) : $signed({{5{w3_mat_real_16[37]}},w3_mat_real_16}); // @[Conditional.scala 39:67 calc6x6.scala 271:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_98 = _T_8 ? $signed(_w3_mat_comp_16_T_8) : $signed({{5{w3_mat_comp_16[37]}},w3_mat_comp_16}); // @[Conditional.scala 39:67 calc6x6.scala 272:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_100 = _T_8 ? $signed({{5{reg2_mat_real_17[19]}},reg2_mat_real_17}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_101 = _T_8 ? $signed(io_weight_real_11) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_11_result = Core_11_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_102 = _T_8 ? $signed(real_11_result) : $signed({{5{w3_mat_real_17[37]}},w3_mat_real_17}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_106 = _T_8 ? $signed(io_weight_comp1_3) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 234:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_107 = _T_8 ? $signed(io_weight_comp2_3) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 235:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_108 = _T_8 ? $signed(io_weight_comp3_3) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 236:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_109 = _T_8 ? $signed({{5{_comp1_3_in_b_T_3[19]}},_comp1_3_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 238:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_110 = _T_8 ? $signed({{5{reg2_mat_real_18[19]}},reg2_mat_real_18}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 239:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_111 = _T_8 ? $signed({{5{reg2_mat_comp_0[19]}},reg2_mat_comp_0}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 240:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_112 = _T_8 ? $signed(_w3_mat_real_18_T_2) : $signed({{5{w3_mat_real_18[37]}},w3_mat_real_18}); // @[Conditional.scala 39:67 calc6x6.scala 241:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_113 = _T_8 ? $signed(_w3_mat_comp_18_T_5) : $signed({{5{w3_mat_comp_18[37]}},w3_mat_comp_18}); // @[Conditional.scala 39:67 calc6x6.scala 242:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_117 = _T_8 ? $signed(io_weight_comp1_4) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 234:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_118 = _T_8 ? $signed(io_weight_comp2_4) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 235:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_119 = _T_8 ? $signed(io_weight_comp3_4) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 236:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_120 = _T_8 ? $signed({{5{_comp1_4_in_b_T_3[19]}},_comp1_4_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 238:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_121 = _T_8 ? $signed({{5{reg2_mat_real_19[19]}},reg2_mat_real_19}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 239:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_122 = _T_8 ? $signed({{5{reg2_mat_comp_1[19]}},reg2_mat_comp_1}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 240:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_123 = _T_8 ? $signed(_w3_mat_real_19_T_2) : $signed({{5{w3_mat_real_19[37]}},w3_mat_real_19}); // @[Conditional.scala 39:67 calc6x6.scala 241:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_124 = _T_8 ? $signed(_w3_mat_comp_19_T_5) : $signed({{5{w3_mat_comp_19[37]}},w3_mat_comp_19}); // @[Conditional.scala 39:67 calc6x6.scala 242:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_128 = _T_8 ? $signed(io_weight_comp1_5) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 234:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_129 = _T_8 ? $signed(io_weight_comp2_5) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 235:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_130 = _T_8 ? $signed(io_weight_comp3_5) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 236:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_131 = _T_8 ? $signed({{5{_comp1_5_in_b_T_3[19]}},_comp1_5_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 238:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_132 = _T_8 ? $signed({{5{reg2_mat_real_20[19]}},reg2_mat_real_20}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 239:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_133 = _T_8 ? $signed({{5{reg2_mat_comp_2[19]}},reg2_mat_comp_2}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 240:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_134 = _T_8 ? $signed(_w3_mat_real_20_T_2) : $signed({{5{w3_mat_real_20[37]}},w3_mat_real_20}); // @[Conditional.scala 39:67 calc6x6.scala 241:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_135 = _T_8 ? $signed(_w3_mat_comp_20_T_5) : $signed({{5{w3_mat_comp_20[37]}},w3_mat_comp_20}); // @[Conditional.scala 39:67 calc6x6.scala 242:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_139 = _T_8 ? $signed(io_weight_comp1_6) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 234:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_140 = _T_8 ? $signed(io_weight_comp2_6) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 235:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_141 = _T_8 ? $signed(io_weight_comp3_6) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 236:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_142 = _T_8 ? $signed({{5{_comp1_6_in_b_T_3[19]}},_comp1_6_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 238:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_143 = _T_8 ? $signed({{5{reg2_mat_real_21[19]}},reg2_mat_real_21}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 239:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_144 = _T_8 ? $signed({{5{reg2_mat_comp_3[19]}},reg2_mat_comp_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 240:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_145 = _T_8 ? $signed(_w3_mat_real_21_T_2) : $signed({{5{w3_mat_real_21[37]}},w3_mat_real_21}); // @[Conditional.scala 39:67 calc6x6.scala 241:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_146 = _T_8 ? $signed(_w3_mat_comp_21_T_5) : $signed({{5{w3_mat_comp_21[37]}},w3_mat_comp_21}); // @[Conditional.scala 39:67 calc6x6.scala 242:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_150 = _T_8 ? $signed(io_weight_comp1_7) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 234:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_151 = _T_8 ? $signed(io_weight_comp2_7) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 235:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_152 = _T_8 ? $signed(io_weight_comp3_7) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 236:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_153 = _T_8 ? $signed({{5{_comp1_7_in_b_T_3[19]}},_comp1_7_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 238:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_154 = _T_8 ? $signed({{5{reg2_mat_real_22[19]}},reg2_mat_real_22}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 239:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_155 = _T_8 ? $signed({{5{reg2_mat_comp_4[19]}},reg2_mat_comp_4}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 240:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_156 = _T_8 ? $signed(_w3_mat_real_22_T_2) : $signed({{5{w3_mat_real_22[37]}},w3_mat_real_22}); // @[Conditional.scala 39:67 calc6x6.scala 241:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_157 = _T_8 ? $signed(_w3_mat_comp_22_T_5) : $signed({{5{w3_mat_comp_22[37]}},w3_mat_comp_22}); // @[Conditional.scala 39:67 calc6x6.scala 242:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_161 = _T_8 ? $signed(io_weight_comp1_8) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 234:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_162 = _T_8 ? $signed(io_weight_comp2_8) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 235:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_163 = _T_8 ? $signed(io_weight_comp3_8) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 236:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_164 = _T_8 ? $signed({{5{_comp1_8_in_b_T_3[19]}},_comp1_8_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 238:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_165 = _T_8 ? $signed({{5{reg2_mat_real_23[19]}},reg2_mat_real_23}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 239:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_166 = _T_8 ? $signed({{5{reg2_mat_comp_5[19]}},reg2_mat_comp_5}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 240:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_167 = _T_8 ? $signed(_w3_mat_real_23_T_2) : $signed({{5{w3_mat_real_23[37]}},w3_mat_real_23}); // @[Conditional.scala 39:67 calc6x6.scala 241:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_168 = _T_8 ? $signed(_w3_mat_comp_23_T_5) : $signed({{5{w3_mat_comp_23[37]}},w3_mat_comp_23}); // @[Conditional.scala 39:67 calc6x6.scala 242:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_169 = _T_8 ? $signed(_w3_mat_real_18_T_2) : $signed({{5{w3_mat_real_24[37]}},w3_mat_real_24}); // @[Conditional.scala 39:67 calc6x6.scala 249:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_170 = _T_8 ? $signed(_w3_mat_comp_24_T_8) : $signed({{5{w3_mat_comp_24[37]}},w3_mat_comp_24}); // @[Conditional.scala 39:67 calc6x6.scala 250:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_171 = _T_8 ? $signed(_w3_mat_real_19_T_2) : $signed({{5{w3_mat_real_25[37]}},w3_mat_real_25}); // @[Conditional.scala 39:67 calc6x6.scala 249:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_172 = _T_8 ? $signed(_w3_mat_comp_25_T_8) : $signed({{5{w3_mat_comp_25[37]}},w3_mat_comp_25}); // @[Conditional.scala 39:67 calc6x6.scala 250:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_173 = _T_8 ? $signed(_w3_mat_real_20_T_2) : $signed({{5{w3_mat_real_26[37]}},w3_mat_real_26}); // @[Conditional.scala 39:67 calc6x6.scala 249:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_174 = _T_8 ? $signed(_w3_mat_comp_26_T_8) : $signed({{5{w3_mat_comp_26[37]}},w3_mat_comp_26}); // @[Conditional.scala 39:67 calc6x6.scala 250:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_175 = _T_8 ? $signed(_w3_mat_real_22_T_2) : $signed({{5{w3_mat_real_27[37]}},w3_mat_real_27}); // @[Conditional.scala 39:67 calc6x6.scala 249:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_176 = _T_8 ? $signed(_w3_mat_comp_27_T_8) : $signed({{5{w3_mat_comp_27[37]}},w3_mat_comp_27}); // @[Conditional.scala 39:67 calc6x6.scala 250:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_177 = _T_8 ? $signed(_w3_mat_real_21_T_2) : $signed({{5{w3_mat_real_28[37]}},w3_mat_real_28}); // @[Conditional.scala 39:67 calc6x6.scala 249:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_178 = _T_8 ? $signed(_w3_mat_comp_28_T_8) : $signed({{5{w3_mat_comp_28[37]}},w3_mat_comp_28}); // @[Conditional.scala 39:67 calc6x6.scala 250:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_179 = _T_8 ? $signed(_w3_mat_real_23_T_2) : $signed({{5{w3_mat_real_29[37]}},w3_mat_real_29}); // @[Conditional.scala 39:67 calc6x6.scala 249:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_180 = _T_8 ? $signed(_w3_mat_comp_29_T_8) : $signed({{5{w3_mat_comp_29[37]}},w3_mat_comp_29}); // @[Conditional.scala 39:67 calc6x6.scala 250:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_182 = _T_8 ? $signed({{5{reg2_mat_real_30[19]}},reg2_mat_real_30}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_183 = _T_8 ? $signed(io_weight_real_12) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_12_result = Core_12_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_184 = _T_8 ? $signed(real_12_result) : $signed({{5{w3_mat_real_30[37]}},w3_mat_real_30}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_186 = _T_8 ? $signed({{5{reg2_mat_real_31[19]}},reg2_mat_real_31}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_187 = _T_8 ? $signed(io_weight_real_13) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_13_result = Core_13_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_188 = _T_8 ? $signed(real_13_result) : $signed({{5{w3_mat_real_31[37]}},w3_mat_real_31}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_190 = _T_8 ? $signed({{5{reg2_mat_real_32[19]}},reg2_mat_real_32}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_191 = _T_8 ? $signed(io_weight_real_14) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_14_result = Core_14_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_192 = _T_8 ? $signed(real_14_result) : $signed({{5{w3_mat_real_32[37]}},w3_mat_real_32}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire [17:0] _GEN_196 = _T_8 ? $signed(io_weight_comp1_9) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 257:38 calc6x6.scala 78:22]
  wire [17:0] _GEN_197 = _T_8 ? $signed(io_weight_comp2_9) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 258:38 calc6x6.scala 81:22]
  wire [17:0] _GEN_198 = _T_8 ? $signed(io_weight_comp3_9) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 259:38 calc6x6.scala 84:22]
  wire [24:0] _GEN_199 = _T_8 ? $signed({{5{_comp1_9_in_b_T_3[19]}},_comp1_9_in_b_T_3}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 261:39 calc6x6.scala 79:23]
  wire [24:0] _GEN_200 = _T_8 ? $signed({{5{reg2_mat_real_33[19]}},reg2_mat_real_33}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 262:39 calc6x6.scala 82:23]
  wire [24:0] _GEN_201 = _T_8 ? $signed({{5{reg2_mat_comp_9[19]}},reg2_mat_comp_9}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 263:39 calc6x6.scala 85:23]
  wire [42:0] _GEN_202 = _T_8 ? $signed(_w3_mat_real_33_T_2) : $signed({{5{w3_mat_real_33[37]}},w3_mat_real_33}); // @[Conditional.scala 39:67 calc6x6.scala 264:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_203 = _T_8 ? $signed(_w3_mat_comp_33_T_5) : $signed({{5{w3_mat_comp_33[37]}},w3_mat_comp_33}); // @[Conditional.scala 39:67 calc6x6.scala 265:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_204 = _T_8 ? $signed(_w3_mat_real_33_T_2) : $signed({{5{w3_mat_real_34[37]}},w3_mat_real_34}); // @[Conditional.scala 39:67 calc6x6.scala 271:47 calc6x6.scala 93:21]
  wire [42:0] _GEN_205 = _T_8 ? $signed(_w3_mat_comp_34_T_8) : $signed({{5{w3_mat_comp_34[37]}},w3_mat_comp_34}); // @[Conditional.scala 39:67 calc6x6.scala 272:47 calc6x6.scala 93:21]
  wire [24:0] _GEN_207 = _T_8 ? $signed({{5{reg2_mat_real_35[19]}},reg2_mat_real_35}) : $signed(25'sh0); // @[Conditional.scala 39:67 calc6x6.scala 225:38 calc6x6.scala 68:22]
  wire [17:0] _GEN_208 = _T_8 ? $signed(io_weight_real_15) : $signed(18'sh0); // @[Conditional.scala 39:67 calc6x6.scala 226:37 calc6x6.scala 67:21]
  wire [42:0] real_15_result = Core_15_io_result; // @[calc6x6.scala 64:23 calc6x6.scala 64:23]
  wire [42:0] _GEN_209 = _T_8 ? $signed(real_15_result) : $signed({{5{w3_mat_real_35[37]}},w3_mat_real_35}); // @[Conditional.scala 39:67 calc6x6.scala 227:47 calc6x6.scala 93:21]
  wire  _GEN_210 = _T_5 | _T_8; // @[Conditional.scala 39:67 calc6x6.scala 195:30]
  wire [24:0] _GEN_211 = _T_5 ? $signed({{9{io_input_mat_0[15]}},io_input_mat_0}) : $signed(_GEN_17); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_212 = _T_5 ? $signed(io_weight_real_0) : $signed(_GEN_18); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_213 = _T_5 ? $signed(real_0_result) : $signed({{5{_GEN_0[37]}},_GEN_0}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_215 = _T_5 ? $signed({{9{io_input_mat_1[15]}},io_input_mat_1}) : $signed(_GEN_21); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_216 = _T_5 ? $signed(io_weight_real_1) : $signed(_GEN_22); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_217 = _T_5 ? $signed(real_1_result) : $signed({{5{_GEN_1[37]}},_GEN_1}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_219 = _T_5 ? $signed({{9{io_input_mat_2[15]}},io_input_mat_2}) : $signed(_GEN_25); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_220 = _T_5 ? $signed(io_weight_real_2) : $signed(_GEN_26); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_221 = _T_5 ? $signed(real_2_result) : $signed({{5{_GEN_2[37]}},_GEN_2}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_223 = _T_5 ? $signed({{9{io_input_mat_3[15]}},io_input_mat_3}) : $signed(_GEN_42); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_224 = _T_5 ? $signed(io_weight_real_3) : $signed(_GEN_43); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_225 = _T_5 ? $signed(real_3_result) : $signed({{5{_GEN_3[37]}},_GEN_3}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_227 = _T_5 ? $signed({{9{io_input_mat_4[15]}},io_input_mat_4}) : $signed(_GEN_46); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_228 = _T_5 ? $signed(io_weight_real_4) : $signed(_GEN_47); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_229 = _T_5 ? $signed(real_4_result) : $signed({{5{_GEN_4[37]}},_GEN_4}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_231 = _T_5 ? $signed({{9{io_input_mat_5[15]}},io_input_mat_5}) : $signed(_GEN_50); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_232 = _T_5 ? $signed(io_weight_real_5) : $signed(_GEN_51); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_233 = _T_5 ? $signed(real_5_result) : $signed({{5{_GEN_5[37]}},_GEN_5}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_235 = _T_5 ? $signed({{9{io_input_mat_6[15]}},io_input_mat_6}) : $signed(_GEN_54); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_236 = _T_5 ? $signed(io_weight_real_6) : $signed(_GEN_55); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_237 = _T_5 ? $signed(real_6_result) : $signed({{5{_GEN_6[37]}},_GEN_6}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_239 = _T_5 ? $signed({{9{io_input_mat_7[15]}},io_input_mat_7}) : $signed(_GEN_71); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_240 = _T_5 ? $signed(io_weight_real_7) : $signed(_GEN_72); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_241 = _T_5 ? $signed(real_7_result) : $signed({{5{_GEN_7[37]}},_GEN_7}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_243 = _T_5 ? $signed({{9{io_input_mat_8[15]}},io_input_mat_8}) : $signed(_GEN_75); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_244 = _T_5 ? $signed(io_weight_real_8) : $signed(_GEN_76); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_245 = _T_5 ? $signed(real_8_result) : $signed({{5{_GEN_8[37]}},_GEN_8}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_247 = _T_5 ? $signed({{9{io_input_mat_9[15]}},io_input_mat_9}) : $signed(_GEN_79); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_248 = _T_5 ? $signed(io_weight_real_9) : $signed(_GEN_80); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_249 = _T_5 ? $signed(real_9_result) : $signed({{5{_GEN_9[37]}},_GEN_9}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_251 = _T_5 ? $signed({{9{io_input_mat_10[15]}},io_input_mat_10}) : $signed(_GEN_83); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_252 = _T_5 ? $signed(io_weight_real_10) : $signed(_GEN_84); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_253 = _T_5 ? $signed(real_10_result) : $signed({{5{_GEN_10[37]}},_GEN_10}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_255 = _T_5 ? $signed({{9{io_input_mat_11[15]}},io_input_mat_11}) : $signed(_GEN_100); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_256 = _T_5 ? $signed(io_weight_real_11) : $signed(_GEN_101); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_257 = _T_5 ? $signed(real_11_result) : $signed({{5{_GEN_11[37]}},_GEN_11}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_259 = _T_5 ? $signed({{9{io_input_mat_12[15]}},io_input_mat_12}) : $signed(_GEN_182); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_260 = _T_5 ? $signed(io_weight_real_12) : $signed(_GEN_183); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_261 = _T_5 ? $signed(real_12_result) : $signed({{5{_GEN_12[37]}},_GEN_12}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_263 = _T_5 ? $signed({{9{io_input_mat_13[15]}},io_input_mat_13}) : $signed(_GEN_186); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_264 = _T_5 ? $signed(io_weight_real_13) : $signed(_GEN_187); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_265 = _T_5 ? $signed(real_13_result) : $signed({{5{_GEN_13[37]}},_GEN_13}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_267 = _T_5 ? $signed({{9{io_input_mat_14[15]}},io_input_mat_14}) : $signed(_GEN_190); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_268 = _T_5 ? $signed(io_weight_real_14) : $signed(_GEN_191); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_269 = _T_5 ? $signed(real_14_result) : $signed({{5{_GEN_14[37]}},_GEN_14}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire [24:0] _GEN_271 = _T_5 ? $signed({{9{io_input_mat_15[15]}},io_input_mat_15}) : $signed(_GEN_207); // @[Conditional.scala 39:67 calc6x6.scala 196:30]
  wire [17:0] _GEN_272 = _T_5 ? $signed(io_weight_real_15) : $signed(_GEN_208); // @[Conditional.scala 39:67 calc6x6.scala 197:29]
  wire [42:0] _GEN_273 = _T_5 ? $signed(real_15_result) : $signed({{5{_GEN_15[37]}},_GEN_15}); // @[Conditional.scala 39:67 calc6x6.scala 198:34]
  wire  _GEN_274 = _T_5 ? io_valid_in : valid_reg_3; // @[Conditional.scala 39:67 calc6x6.scala 201:25 calc6x6.scala 180:18]
  wire [42:0] _GEN_275 = _T_5 ? $signed({{5{w3_mat_real_0[37]}},w3_mat_real_0}) : $signed(_GEN_19); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_276 = _T_5 ? $signed({{5{w3_mat_real_1[37]}},w3_mat_real_1}) : $signed(_GEN_23); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_277 = _T_5 ? $signed({{5{w3_mat_real_2[37]}},w3_mat_real_2}) : $signed(_GEN_27); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire  _GEN_278 = _T_5 ? 1'h0 : _T_8; // @[Conditional.scala 39:67 calc6x6.scala 77:23]
  wire [17:0] _GEN_281 = _T_5 ? $signed(18'sh0) : $signed(_GEN_31); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_282 = _T_5 ? $signed(18'sh0) : $signed(_GEN_32); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_283 = _T_5 ? $signed(18'sh0) : $signed(_GEN_33); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_284 = _T_5 ? $signed(25'sh0) : $signed(_GEN_34); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_285 = _T_5 ? $signed(25'sh0) : $signed(_GEN_35); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_286 = _T_5 ? $signed(25'sh0) : $signed(_GEN_36); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_287 = _T_5 ? $signed({{5{w3_mat_real_3[37]}},w3_mat_real_3}) : $signed(_GEN_37); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_288 = _T_5 ? $signed({{5{w3_mat_comp_3[37]}},w3_mat_comp_3}) : $signed(_GEN_38); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_289 = _T_5 ? $signed({{5{w3_mat_real_4[37]}},w3_mat_real_4}) : $signed(_GEN_39); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_290 = _T_5 ? $signed({{5{w3_mat_comp_4[37]}},w3_mat_comp_4}) : $signed(_GEN_40); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_291 = _T_5 ? $signed({{5{w3_mat_real_5[37]}},w3_mat_real_5}) : $signed(_GEN_44); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_292 = _T_5 ? $signed({{5{w3_mat_real_6[37]}},w3_mat_real_6}) : $signed(_GEN_48); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_293 = _T_5 ? $signed({{5{w3_mat_real_7[37]}},w3_mat_real_7}) : $signed(_GEN_52); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_294 = _T_5 ? $signed({{5{w3_mat_real_8[37]}},w3_mat_real_8}) : $signed(_GEN_56); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_298 = _T_5 ? $signed(18'sh0) : $signed(_GEN_60); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_299 = _T_5 ? $signed(18'sh0) : $signed(_GEN_61); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_300 = _T_5 ? $signed(18'sh0) : $signed(_GEN_62); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_301 = _T_5 ? $signed(25'sh0) : $signed(_GEN_63); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_302 = _T_5 ? $signed(25'sh0) : $signed(_GEN_64); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_303 = _T_5 ? $signed(25'sh0) : $signed(_GEN_65); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_304 = _T_5 ? $signed({{5{w3_mat_real_9[37]}},w3_mat_real_9}) : $signed(_GEN_66); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_305 = _T_5 ? $signed({{5{w3_mat_comp_9[37]}},w3_mat_comp_9}) : $signed(_GEN_67); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_306 = _T_5 ? $signed({{5{w3_mat_real_10[37]}},w3_mat_real_10}) : $signed(_GEN_68); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_307 = _T_5 ? $signed({{5{w3_mat_comp_10[37]}},w3_mat_comp_10}) : $signed(_GEN_69); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_308 = _T_5 ? $signed({{5{w3_mat_real_11[37]}},w3_mat_real_11}) : $signed(_GEN_73); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_309 = _T_5 ? $signed({{5{w3_mat_real_12[37]}},w3_mat_real_12}) : $signed(_GEN_77); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_310 = _T_5 ? $signed({{5{w3_mat_real_13[37]}},w3_mat_real_13}) : $signed(_GEN_81); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_311 = _T_5 ? $signed({{5{w3_mat_real_14[37]}},w3_mat_real_14}) : $signed(_GEN_85); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_315 = _T_5 ? $signed(18'sh0) : $signed(_GEN_89); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_316 = _T_5 ? $signed(18'sh0) : $signed(_GEN_90); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_317 = _T_5 ? $signed(18'sh0) : $signed(_GEN_91); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_318 = _T_5 ? $signed(25'sh0) : $signed(_GEN_92); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_319 = _T_5 ? $signed(25'sh0) : $signed(_GEN_93); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_320 = _T_5 ? $signed(25'sh0) : $signed(_GEN_94); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_321 = _T_5 ? $signed({{5{w3_mat_real_15[37]}},w3_mat_real_15}) : $signed(_GEN_95); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_322 = _T_5 ? $signed({{5{w3_mat_comp_15[37]}},w3_mat_comp_15}) : $signed(_GEN_96); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_323 = _T_5 ? $signed({{5{w3_mat_real_16[37]}},w3_mat_real_16}) : $signed(_GEN_97); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_324 = _T_5 ? $signed({{5{w3_mat_comp_16[37]}},w3_mat_comp_16}) : $signed(_GEN_98); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_325 = _T_5 ? $signed({{5{w3_mat_real_17[37]}},w3_mat_real_17}) : $signed(_GEN_102); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_329 = _T_5 ? $signed(18'sh0) : $signed(_GEN_106); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_330 = _T_5 ? $signed(18'sh0) : $signed(_GEN_107); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_331 = _T_5 ? $signed(18'sh0) : $signed(_GEN_108); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_332 = _T_5 ? $signed(25'sh0) : $signed(_GEN_109); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_333 = _T_5 ? $signed(25'sh0) : $signed(_GEN_110); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_334 = _T_5 ? $signed(25'sh0) : $signed(_GEN_111); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_335 = _T_5 ? $signed({{5{w3_mat_real_18[37]}},w3_mat_real_18}) : $signed(_GEN_112); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_336 = _T_5 ? $signed({{5{w3_mat_comp_18[37]}},w3_mat_comp_18}) : $signed(_GEN_113); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_340 = _T_5 ? $signed(18'sh0) : $signed(_GEN_117); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_341 = _T_5 ? $signed(18'sh0) : $signed(_GEN_118); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_342 = _T_5 ? $signed(18'sh0) : $signed(_GEN_119); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_343 = _T_5 ? $signed(25'sh0) : $signed(_GEN_120); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_344 = _T_5 ? $signed(25'sh0) : $signed(_GEN_121); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_345 = _T_5 ? $signed(25'sh0) : $signed(_GEN_122); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_346 = _T_5 ? $signed({{5{w3_mat_real_19[37]}},w3_mat_real_19}) : $signed(_GEN_123); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_347 = _T_5 ? $signed({{5{w3_mat_comp_19[37]}},w3_mat_comp_19}) : $signed(_GEN_124); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_351 = _T_5 ? $signed(18'sh0) : $signed(_GEN_128); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_352 = _T_5 ? $signed(18'sh0) : $signed(_GEN_129); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_353 = _T_5 ? $signed(18'sh0) : $signed(_GEN_130); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_354 = _T_5 ? $signed(25'sh0) : $signed(_GEN_131); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_355 = _T_5 ? $signed(25'sh0) : $signed(_GEN_132); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_356 = _T_5 ? $signed(25'sh0) : $signed(_GEN_133); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_357 = _T_5 ? $signed({{5{w3_mat_real_20[37]}},w3_mat_real_20}) : $signed(_GEN_134); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_358 = _T_5 ? $signed({{5{w3_mat_comp_20[37]}},w3_mat_comp_20}) : $signed(_GEN_135); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_362 = _T_5 ? $signed(18'sh0) : $signed(_GEN_139); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_363 = _T_5 ? $signed(18'sh0) : $signed(_GEN_140); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_364 = _T_5 ? $signed(18'sh0) : $signed(_GEN_141); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_365 = _T_5 ? $signed(25'sh0) : $signed(_GEN_142); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_366 = _T_5 ? $signed(25'sh0) : $signed(_GEN_143); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_367 = _T_5 ? $signed(25'sh0) : $signed(_GEN_144); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_368 = _T_5 ? $signed({{5{w3_mat_real_21[37]}},w3_mat_real_21}) : $signed(_GEN_145); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_369 = _T_5 ? $signed({{5{w3_mat_comp_21[37]}},w3_mat_comp_21}) : $signed(_GEN_146); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_373 = _T_5 ? $signed(18'sh0) : $signed(_GEN_150); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_374 = _T_5 ? $signed(18'sh0) : $signed(_GEN_151); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_375 = _T_5 ? $signed(18'sh0) : $signed(_GEN_152); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_376 = _T_5 ? $signed(25'sh0) : $signed(_GEN_153); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_377 = _T_5 ? $signed(25'sh0) : $signed(_GEN_154); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_378 = _T_5 ? $signed(25'sh0) : $signed(_GEN_155); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_379 = _T_5 ? $signed({{5{w3_mat_real_22[37]}},w3_mat_real_22}) : $signed(_GEN_156); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_380 = _T_5 ? $signed({{5{w3_mat_comp_22[37]}},w3_mat_comp_22}) : $signed(_GEN_157); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_384 = _T_5 ? $signed(18'sh0) : $signed(_GEN_161); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_385 = _T_5 ? $signed(18'sh0) : $signed(_GEN_162); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_386 = _T_5 ? $signed(18'sh0) : $signed(_GEN_163); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_387 = _T_5 ? $signed(25'sh0) : $signed(_GEN_164); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_388 = _T_5 ? $signed(25'sh0) : $signed(_GEN_165); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_389 = _T_5 ? $signed(25'sh0) : $signed(_GEN_166); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_390 = _T_5 ? $signed({{5{w3_mat_real_23[37]}},w3_mat_real_23}) : $signed(_GEN_167); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_391 = _T_5 ? $signed({{5{w3_mat_comp_23[37]}},w3_mat_comp_23}) : $signed(_GEN_168); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_392 = _T_5 ? $signed({{5{w3_mat_real_24[37]}},w3_mat_real_24}) : $signed(_GEN_169); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_393 = _T_5 ? $signed({{5{w3_mat_comp_24[37]}},w3_mat_comp_24}) : $signed(_GEN_170); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_394 = _T_5 ? $signed({{5{w3_mat_real_25[37]}},w3_mat_real_25}) : $signed(_GEN_171); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_395 = _T_5 ? $signed({{5{w3_mat_comp_25[37]}},w3_mat_comp_25}) : $signed(_GEN_172); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_396 = _T_5 ? $signed({{5{w3_mat_real_26[37]}},w3_mat_real_26}) : $signed(_GEN_173); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_397 = _T_5 ? $signed({{5{w3_mat_comp_26[37]}},w3_mat_comp_26}) : $signed(_GEN_174); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_398 = _T_5 ? $signed({{5{w3_mat_real_27[37]}},w3_mat_real_27}) : $signed(_GEN_175); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_399 = _T_5 ? $signed({{5{w3_mat_comp_27[37]}},w3_mat_comp_27}) : $signed(_GEN_176); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_400 = _T_5 ? $signed({{5{w3_mat_real_28[37]}},w3_mat_real_28}) : $signed(_GEN_177); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_401 = _T_5 ? $signed({{5{w3_mat_comp_28[37]}},w3_mat_comp_28}) : $signed(_GEN_178); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_402 = _T_5 ? $signed({{5{w3_mat_real_29[37]}},w3_mat_real_29}) : $signed(_GEN_179); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_403 = _T_5 ? $signed({{5{w3_mat_comp_29[37]}},w3_mat_comp_29}) : $signed(_GEN_180); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_404 = _T_5 ? $signed({{5{w3_mat_real_30[37]}},w3_mat_real_30}) : $signed(_GEN_184); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_405 = _T_5 ? $signed({{5{w3_mat_real_31[37]}},w3_mat_real_31}) : $signed(_GEN_188); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_406 = _T_5 ? $signed({{5{w3_mat_real_32[37]}},w3_mat_real_32}) : $signed(_GEN_192); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [17:0] _GEN_410 = _T_5 ? $signed(18'sh0) : $signed(_GEN_196); // @[Conditional.scala 39:67 calc6x6.scala 78:22]
  wire [17:0] _GEN_411 = _T_5 ? $signed(18'sh0) : $signed(_GEN_197); // @[Conditional.scala 39:67 calc6x6.scala 81:22]
  wire [17:0] _GEN_412 = _T_5 ? $signed(18'sh0) : $signed(_GEN_198); // @[Conditional.scala 39:67 calc6x6.scala 84:22]
  wire [24:0] _GEN_413 = _T_5 ? $signed(25'sh0) : $signed(_GEN_199); // @[Conditional.scala 39:67 calc6x6.scala 79:23]
  wire [24:0] _GEN_414 = _T_5 ? $signed(25'sh0) : $signed(_GEN_200); // @[Conditional.scala 39:67 calc6x6.scala 82:23]
  wire [24:0] _GEN_415 = _T_5 ? $signed(25'sh0) : $signed(_GEN_201); // @[Conditional.scala 39:67 calc6x6.scala 85:23]
  wire [42:0] _GEN_416 = _T_5 ? $signed({{5{w3_mat_real_33[37]}},w3_mat_real_33}) : $signed(_GEN_202); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_417 = _T_5 ? $signed({{5{w3_mat_comp_33[37]}},w3_mat_comp_33}) : $signed(_GEN_203); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_418 = _T_5 ? $signed({{5{w3_mat_real_34[37]}},w3_mat_real_34}) : $signed(_GEN_204); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_419 = _T_5 ? $signed({{5{w3_mat_comp_34[37]}},w3_mat_comp_34}) : $signed(_GEN_205); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_420 = _T_5 ? $signed({{5{w3_mat_real_35[37]}},w3_mat_real_35}) : $signed(_GEN_209); // @[Conditional.scala 39:67 calc6x6.scala 93:21]
  wire [42:0] _GEN_423 = _T_2 ? $signed(real_0_result) : $signed(_GEN_213); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_426 = _T_2 ? $signed(real_1_result) : $signed(_GEN_217); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_429 = _T_2 ? $signed(real_2_result) : $signed(_GEN_221); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_432 = _T_2 ? $signed(real_3_result) : $signed(_GEN_225); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_435 = _T_2 ? $signed(real_4_result) : $signed(_GEN_229); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_438 = _T_2 ? $signed(real_5_result) : $signed(_GEN_233); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_441 = _T_2 ? $signed(real_6_result) : $signed(_GEN_237); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_444 = _T_2 ? $signed(real_7_result) : $signed(_GEN_241); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_447 = _T_2 ? $signed(real_8_result) : $signed(_GEN_245); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_450 = _T_2 ? $signed(real_9_result) : $signed(_GEN_249); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_453 = _T_2 ? $signed(real_10_result) : $signed(_GEN_253); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_456 = _T_2 ? $signed(real_11_result) : $signed(_GEN_257); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_459 = _T_2 ? $signed(real_12_result) : $signed(_GEN_261); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_462 = _T_2 ? $signed(real_13_result) : $signed(_GEN_265); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_465 = _T_2 ? $signed(real_14_result) : $signed(_GEN_269); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_468 = _T_2 ? $signed(real_15_result) : $signed(_GEN_273); // @[Conditional.scala 40:58 calc6x6.scala 187:34]
  wire [42:0] _GEN_486 = _T_2 ? $signed({{5{w3_mat_real_0[37]}},w3_mat_real_0}) : $signed(_GEN_275); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_487 = _T_2 ? $signed({{5{w3_mat_real_1[37]}},w3_mat_real_1}) : $signed(_GEN_276); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_488 = _T_2 ? $signed({{5{w3_mat_real_2[37]}},w3_mat_real_2}) : $signed(_GEN_277); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_498 = _T_2 ? $signed({{5{w3_mat_real_3[37]}},w3_mat_real_3}) : $signed(_GEN_287); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_499 = _T_2 ? $signed({{5{w3_mat_comp_3[37]}},w3_mat_comp_3}) : $signed(_GEN_288); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_500 = _T_2 ? $signed({{5{w3_mat_real_4[37]}},w3_mat_real_4}) : $signed(_GEN_289); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_501 = _T_2 ? $signed({{5{w3_mat_comp_4[37]}},w3_mat_comp_4}) : $signed(_GEN_290); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_502 = _T_2 ? $signed({{5{w3_mat_real_5[37]}},w3_mat_real_5}) : $signed(_GEN_291); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_503 = _T_2 ? $signed({{5{w3_mat_real_6[37]}},w3_mat_real_6}) : $signed(_GEN_292); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_504 = _T_2 ? $signed({{5{w3_mat_real_7[37]}},w3_mat_real_7}) : $signed(_GEN_293); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_505 = _T_2 ? $signed({{5{w3_mat_real_8[37]}},w3_mat_real_8}) : $signed(_GEN_294); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_515 = _T_2 ? $signed({{5{w3_mat_real_9[37]}},w3_mat_real_9}) : $signed(_GEN_304); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_516 = _T_2 ? $signed({{5{w3_mat_comp_9[37]}},w3_mat_comp_9}) : $signed(_GEN_305); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_517 = _T_2 ? $signed({{5{w3_mat_real_10[37]}},w3_mat_real_10}) : $signed(_GEN_306); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_518 = _T_2 ? $signed({{5{w3_mat_comp_10[37]}},w3_mat_comp_10}) : $signed(_GEN_307); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_519 = _T_2 ? $signed({{5{w3_mat_real_11[37]}},w3_mat_real_11}) : $signed(_GEN_308); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_520 = _T_2 ? $signed({{5{w3_mat_real_12[37]}},w3_mat_real_12}) : $signed(_GEN_309); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_521 = _T_2 ? $signed({{5{w3_mat_real_13[37]}},w3_mat_real_13}) : $signed(_GEN_310); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_522 = _T_2 ? $signed({{5{w3_mat_real_14[37]}},w3_mat_real_14}) : $signed(_GEN_311); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_532 = _T_2 ? $signed({{5{w3_mat_real_15[37]}},w3_mat_real_15}) : $signed(_GEN_321); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_533 = _T_2 ? $signed({{5{w3_mat_comp_15[37]}},w3_mat_comp_15}) : $signed(_GEN_322); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_534 = _T_2 ? $signed({{5{w3_mat_real_16[37]}},w3_mat_real_16}) : $signed(_GEN_323); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_535 = _T_2 ? $signed({{5{w3_mat_comp_16[37]}},w3_mat_comp_16}) : $signed(_GEN_324); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_536 = _T_2 ? $signed({{5{w3_mat_real_17[37]}},w3_mat_real_17}) : $signed(_GEN_325); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_546 = _T_2 ? $signed({{5{w3_mat_real_18[37]}},w3_mat_real_18}) : $signed(_GEN_335); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_547 = _T_2 ? $signed({{5{w3_mat_comp_18[37]}},w3_mat_comp_18}) : $signed(_GEN_336); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_557 = _T_2 ? $signed({{5{w3_mat_real_19[37]}},w3_mat_real_19}) : $signed(_GEN_346); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_558 = _T_2 ? $signed({{5{w3_mat_comp_19[37]}},w3_mat_comp_19}) : $signed(_GEN_347); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_568 = _T_2 ? $signed({{5{w3_mat_real_20[37]}},w3_mat_real_20}) : $signed(_GEN_357); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_569 = _T_2 ? $signed({{5{w3_mat_comp_20[37]}},w3_mat_comp_20}) : $signed(_GEN_358); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_579 = _T_2 ? $signed({{5{w3_mat_real_21[37]}},w3_mat_real_21}) : $signed(_GEN_368); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_580 = _T_2 ? $signed({{5{w3_mat_comp_21[37]}},w3_mat_comp_21}) : $signed(_GEN_369); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_590 = _T_2 ? $signed({{5{w3_mat_real_22[37]}},w3_mat_real_22}) : $signed(_GEN_379); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_591 = _T_2 ? $signed({{5{w3_mat_comp_22[37]}},w3_mat_comp_22}) : $signed(_GEN_380); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_601 = _T_2 ? $signed({{5{w3_mat_real_23[37]}},w3_mat_real_23}) : $signed(_GEN_390); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_602 = _T_2 ? $signed({{5{w3_mat_comp_23[37]}},w3_mat_comp_23}) : $signed(_GEN_391); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_603 = _T_2 ? $signed({{5{w3_mat_real_24[37]}},w3_mat_real_24}) : $signed(_GEN_392); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_604 = _T_2 ? $signed({{5{w3_mat_comp_24[37]}},w3_mat_comp_24}) : $signed(_GEN_393); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_605 = _T_2 ? $signed({{5{w3_mat_real_25[37]}},w3_mat_real_25}) : $signed(_GEN_394); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_606 = _T_2 ? $signed({{5{w3_mat_comp_25[37]}},w3_mat_comp_25}) : $signed(_GEN_395); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_607 = _T_2 ? $signed({{5{w3_mat_real_26[37]}},w3_mat_real_26}) : $signed(_GEN_396); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_608 = _T_2 ? $signed({{5{w3_mat_comp_26[37]}},w3_mat_comp_26}) : $signed(_GEN_397); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_609 = _T_2 ? $signed({{5{w3_mat_real_27[37]}},w3_mat_real_27}) : $signed(_GEN_398); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_610 = _T_2 ? $signed({{5{w3_mat_comp_27[37]}},w3_mat_comp_27}) : $signed(_GEN_399); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_611 = _T_2 ? $signed({{5{w3_mat_real_28[37]}},w3_mat_real_28}) : $signed(_GEN_400); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_612 = _T_2 ? $signed({{5{w3_mat_comp_28[37]}},w3_mat_comp_28}) : $signed(_GEN_401); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_613 = _T_2 ? $signed({{5{w3_mat_real_29[37]}},w3_mat_real_29}) : $signed(_GEN_402); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_614 = _T_2 ? $signed({{5{w3_mat_comp_29[37]}},w3_mat_comp_29}) : $signed(_GEN_403); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_615 = _T_2 ? $signed({{5{w3_mat_real_30[37]}},w3_mat_real_30}) : $signed(_GEN_404); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_616 = _T_2 ? $signed({{5{w3_mat_real_31[37]}},w3_mat_real_31}) : $signed(_GEN_405); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_617 = _T_2 ? $signed({{5{w3_mat_real_32[37]}},w3_mat_real_32}) : $signed(_GEN_406); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_627 = _T_2 ? $signed({{5{w3_mat_real_33[37]}},w3_mat_real_33}) : $signed(_GEN_416); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_628 = _T_2 ? $signed({{5{w3_mat_comp_33[37]}},w3_mat_comp_33}) : $signed(_GEN_417); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_629 = _T_2 ? $signed({{5{w3_mat_real_34[37]}},w3_mat_real_34}) : $signed(_GEN_418); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_630 = _T_2 ? $signed({{5{w3_mat_comp_34[37]}},w3_mat_comp_34}) : $signed(_GEN_419); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  wire [42:0] _GEN_631 = _T_2 ? $signed({{5{w3_mat_real_35[37]}},w3_mat_real_35}) : $signed(_GEN_420); // @[Conditional.scala 40:58 calc6x6.scala 93:21]
  Core Core ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_io_w_a),
    .io_in_b(Core_io_in_b),
    .io_flag(Core_io_flag),
    .io_result(Core_io_result)
  );
  Core Core_1 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_1_io_w_a),
    .io_in_b(Core_1_io_in_b),
    .io_flag(Core_1_io_flag),
    .io_result(Core_1_io_result)
  );
  Core Core_2 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_2_io_w_a),
    .io_in_b(Core_2_io_in_b),
    .io_flag(Core_2_io_flag),
    .io_result(Core_2_io_result)
  );
  Core Core_3 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_3_io_w_a),
    .io_in_b(Core_3_io_in_b),
    .io_flag(Core_3_io_flag),
    .io_result(Core_3_io_result)
  );
  Core Core_4 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_4_io_w_a),
    .io_in_b(Core_4_io_in_b),
    .io_flag(Core_4_io_flag),
    .io_result(Core_4_io_result)
  );
  Core Core_5 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_5_io_w_a),
    .io_in_b(Core_5_io_in_b),
    .io_flag(Core_5_io_flag),
    .io_result(Core_5_io_result)
  );
  Core Core_6 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_6_io_w_a),
    .io_in_b(Core_6_io_in_b),
    .io_flag(Core_6_io_flag),
    .io_result(Core_6_io_result)
  );
  Core Core_7 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_7_io_w_a),
    .io_in_b(Core_7_io_in_b),
    .io_flag(Core_7_io_flag),
    .io_result(Core_7_io_result)
  );
  Core Core_8 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_8_io_w_a),
    .io_in_b(Core_8_io_in_b),
    .io_flag(Core_8_io_flag),
    .io_result(Core_8_io_result)
  );
  Core Core_9 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_9_io_w_a),
    .io_in_b(Core_9_io_in_b),
    .io_flag(Core_9_io_flag),
    .io_result(Core_9_io_result)
  );
  Core Core_10 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_10_io_w_a),
    .io_in_b(Core_10_io_in_b),
    .io_flag(Core_10_io_flag),
    .io_result(Core_10_io_result)
  );
  Core Core_11 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_11_io_w_a),
    .io_in_b(Core_11_io_in_b),
    .io_flag(Core_11_io_flag),
    .io_result(Core_11_io_result)
  );
  Core Core_12 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_12_io_w_a),
    .io_in_b(Core_12_io_in_b),
    .io_flag(Core_12_io_flag),
    .io_result(Core_12_io_result)
  );
  Core Core_13 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_13_io_w_a),
    .io_in_b(Core_13_io_in_b),
    .io_flag(Core_13_io_flag),
    .io_result(Core_13_io_result)
  );
  Core Core_14 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_14_io_w_a),
    .io_in_b(Core_14_io_in_b),
    .io_flag(Core_14_io_flag),
    .io_result(Core_14_io_result)
  );
  Core Core_15 ( // @[calc6x6.scala 64:43]
    .io_w_a(Core_15_io_w_a),
    .io_in_b(Core_15_io_in_b),
    .io_flag(Core_15_io_flag),
    .io_result(Core_15_io_result)
  );
  Core Core_16 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_16_io_w_a),
    .io_in_b(Core_16_io_in_b),
    .io_flag(Core_16_io_flag),
    .io_result(Core_16_io_result)
  );
  Core Core_17 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_17_io_w_a),
    .io_in_b(Core_17_io_in_b),
    .io_flag(Core_17_io_flag),
    .io_result(Core_17_io_result)
  );
  Core Core_18 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_18_io_w_a),
    .io_in_b(Core_18_io_in_b),
    .io_flag(Core_18_io_flag),
    .io_result(Core_18_io_result)
  );
  Core Core_19 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_19_io_w_a),
    .io_in_b(Core_19_io_in_b),
    .io_flag(Core_19_io_flag),
    .io_result(Core_19_io_result)
  );
  Core Core_20 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_20_io_w_a),
    .io_in_b(Core_20_io_in_b),
    .io_flag(Core_20_io_flag),
    .io_result(Core_20_io_result)
  );
  Core Core_21 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_21_io_w_a),
    .io_in_b(Core_21_io_in_b),
    .io_flag(Core_21_io_flag),
    .io_result(Core_21_io_result)
  );
  Core Core_22 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_22_io_w_a),
    .io_in_b(Core_22_io_in_b),
    .io_flag(Core_22_io_flag),
    .io_result(Core_22_io_result)
  );
  Core Core_23 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_23_io_w_a),
    .io_in_b(Core_23_io_in_b),
    .io_flag(Core_23_io_flag),
    .io_result(Core_23_io_result)
  );
  Core Core_24 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_24_io_w_a),
    .io_in_b(Core_24_io_in_b),
    .io_flag(Core_24_io_flag),
    .io_result(Core_24_io_result)
  );
  Core Core_25 ( // @[calc6x6.scala 71:44]
    .io_w_a(Core_25_io_w_a),
    .io_in_b(Core_25_io_in_b),
    .io_flag(Core_25_io_flag),
    .io_result(Core_25_io_result)
  );
  Core Core_26 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_26_io_w_a),
    .io_in_b(Core_26_io_in_b),
    .io_flag(Core_26_io_flag),
    .io_result(Core_26_io_result)
  );
  Core Core_27 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_27_io_w_a),
    .io_in_b(Core_27_io_in_b),
    .io_flag(Core_27_io_flag),
    .io_result(Core_27_io_result)
  );
  Core Core_28 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_28_io_w_a),
    .io_in_b(Core_28_io_in_b),
    .io_flag(Core_28_io_flag),
    .io_result(Core_28_io_result)
  );
  Core Core_29 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_29_io_w_a),
    .io_in_b(Core_29_io_in_b),
    .io_flag(Core_29_io_flag),
    .io_result(Core_29_io_result)
  );
  Core Core_30 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_30_io_w_a),
    .io_in_b(Core_30_io_in_b),
    .io_flag(Core_30_io_flag),
    .io_result(Core_30_io_result)
  );
  Core Core_31 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_31_io_w_a),
    .io_in_b(Core_31_io_in_b),
    .io_flag(Core_31_io_flag),
    .io_result(Core_31_io_result)
  );
  Core Core_32 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_32_io_w_a),
    .io_in_b(Core_32_io_in_b),
    .io_flag(Core_32_io_flag),
    .io_result(Core_32_io_result)
  );
  Core Core_33 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_33_io_w_a),
    .io_in_b(Core_33_io_in_b),
    .io_flag(Core_33_io_flag),
    .io_result(Core_33_io_result)
  );
  Core Core_34 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_34_io_w_a),
    .io_in_b(Core_34_io_in_b),
    .io_flag(Core_34_io_flag),
    .io_result(Core_34_io_result)
  );
  Core Core_35 ( // @[calc6x6.scala 72:44]
    .io_w_a(Core_35_io_w_a),
    .io_in_b(Core_35_io_in_b),
    .io_flag(Core_35_io_flag),
    .io_result(Core_35_io_result)
  );
  Core Core_36 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_36_io_w_a),
    .io_in_b(Core_36_io_in_b),
    .io_flag(Core_36_io_flag),
    .io_result(Core_36_io_result)
  );
  Core Core_37 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_37_io_w_a),
    .io_in_b(Core_37_io_in_b),
    .io_flag(Core_37_io_flag),
    .io_result(Core_37_io_result)
  );
  Core Core_38 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_38_io_w_a),
    .io_in_b(Core_38_io_in_b),
    .io_flag(Core_38_io_flag),
    .io_result(Core_38_io_result)
  );
  Core Core_39 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_39_io_w_a),
    .io_in_b(Core_39_io_in_b),
    .io_flag(Core_39_io_flag),
    .io_result(Core_39_io_result)
  );
  Core Core_40 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_40_io_w_a),
    .io_in_b(Core_40_io_in_b),
    .io_flag(Core_40_io_flag),
    .io_result(Core_40_io_result)
  );
  Core Core_41 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_41_io_w_a),
    .io_in_b(Core_41_io_in_b),
    .io_flag(Core_41_io_flag),
    .io_result(Core_41_io_result)
  );
  Core Core_42 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_42_io_w_a),
    .io_in_b(Core_42_io_in_b),
    .io_flag(Core_42_io_flag),
    .io_result(Core_42_io_result)
  );
  Core Core_43 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_43_io_w_a),
    .io_in_b(Core_43_io_in_b),
    .io_flag(Core_43_io_flag),
    .io_result(Core_43_io_result)
  );
  Core Core_44 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_44_io_w_a),
    .io_in_b(Core_44_io_in_b),
    .io_flag(Core_44_io_flag),
    .io_result(Core_44_io_result)
  );
  Core Core_45 ( // @[calc6x6.scala 73:44]
    .io_w_a(Core_45_io_w_a),
    .io_in_b(Core_45_io_in_b),
    .io_flag(Core_45_io_flag),
    .io_result(Core_45_io_result)
  );
  assign io_output_mat_0 = _GEN_423[36:0];
  assign io_output_mat_1 = _GEN_426[36:0];
  assign io_output_mat_2 = _GEN_429[36:0];
  assign io_output_mat_3 = _GEN_432[36:0];
  assign io_output_mat_4 = _GEN_435[36:0];
  assign io_output_mat_5 = _GEN_438[36:0];
  assign io_output_mat_6 = _GEN_441[36:0];
  assign io_output_mat_7 = _GEN_444[36:0];
  assign io_output_mat_8 = _GEN_447[36:0];
  assign io_output_mat_9 = _GEN_450[36:0];
  assign io_output_mat_10 = _GEN_453[36:0];
  assign io_output_mat_11 = _GEN_456[36:0];
  assign io_output_mat_12 = _GEN_459[36:0];
  assign io_output_mat_13 = _GEN_462[36:0];
  assign io_output_mat_14 = _GEN_465[36:0];
  assign io_output_mat_15 = _GEN_468[36:0];
  assign io_valid_out = _T_2 ? io_valid_in : _GEN_274; // @[Conditional.scala 40:58 calc6x6.scala 189:26]
  assign Core_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_212); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_io_in_b = _T_2 ? $signed({{9{io_input_mat_0[15]}},io_input_mat_0}) : $signed(_GEN_211); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_1_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_216); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_1_io_in_b = _T_2 ? $signed({{9{io_input_mat_1[15]}},io_input_mat_1}) : $signed(_GEN_215); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_1_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_2_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_220); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_2_io_in_b = _T_2 ? $signed({{9{io_input_mat_2[15]}},io_input_mat_2}) : $signed(_GEN_219); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_2_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_3_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_224); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_3_io_in_b = _T_2 ? $signed({{9{io_input_mat_3[15]}},io_input_mat_3}) : $signed(_GEN_223); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_3_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_4_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_228); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_4_io_in_b = _T_2 ? $signed({{9{io_input_mat_4[15]}},io_input_mat_4}) : $signed(_GEN_227); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_4_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_5_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_232); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_5_io_in_b = _T_2 ? $signed({{9{io_input_mat_5[15]}},io_input_mat_5}) : $signed(_GEN_231); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_5_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_6_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_236); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_6_io_in_b = _T_2 ? $signed({{9{io_input_mat_6[15]}},io_input_mat_6}) : $signed(_GEN_235); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_6_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_7_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_240); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_7_io_in_b = _T_2 ? $signed({{9{io_input_mat_7[15]}},io_input_mat_7}) : $signed(_GEN_239); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_7_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_8_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_244); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_8_io_in_b = _T_2 ? $signed({{9{io_input_mat_8[15]}},io_input_mat_8}) : $signed(_GEN_243); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_8_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_9_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_248); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_9_io_in_b = _T_2 ? $signed({{9{io_input_mat_9[15]}},io_input_mat_9}) : $signed(_GEN_247); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_9_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_10_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_252); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_10_io_in_b = _T_2 ? $signed({{9{io_input_mat_10[15]}},io_input_mat_10}) : $signed(_GEN_251); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_10_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_11_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_256); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_11_io_in_b = _T_2 ? $signed({{9{io_input_mat_11[15]}},io_input_mat_11}) : $signed(_GEN_255); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_11_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_12_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_260); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_12_io_in_b = _T_2 ? $signed({{9{io_input_mat_12[15]}},io_input_mat_12}) : $signed(_GEN_259); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_12_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_13_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_264); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_13_io_in_b = _T_2 ? $signed({{9{io_input_mat_13[15]}},io_input_mat_13}) : $signed(_GEN_263); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_13_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_14_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_268); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_14_io_in_b = _T_2 ? $signed({{9{io_input_mat_14[15]}},io_input_mat_14}) : $signed(_GEN_267); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_14_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_15_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_272); // @[Conditional.scala 40:58 calc6x6.scala 67:21]
  assign Core_15_io_in_b = _T_2 ? $signed({{9{io_input_mat_15[15]}},io_input_mat_15}) : $signed(_GEN_271); // @[Conditional.scala 40:58 calc6x6.scala 186:30]
  assign Core_15_io_flag = _T_2 ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58 calc6x6.scala 185:30]
  assign Core_16_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_281); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_16_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_284); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_16_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_17_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_298); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_17_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_301); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_17_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_18_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_315); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_18_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_318); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_18_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_19_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_329); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_19_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_332); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_19_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_20_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_340); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_20_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_343); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_20_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_21_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_351); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_21_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_354); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_21_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_22_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_362); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_22_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_365); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_22_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_23_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_373); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_23_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_376); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_23_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_24_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_384); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_24_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_387); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_24_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_25_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_410); // @[Conditional.scala 40:58 calc6x6.scala 78:22]
  assign Core_25_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_413); // @[Conditional.scala 40:58 calc6x6.scala 79:23]
  assign Core_25_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 77:23]
  assign Core_26_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_282); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_26_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_285); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_26_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_27_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_299); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_27_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_302); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_27_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_28_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_316); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_28_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_319); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_28_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_29_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_330); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_29_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_333); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_29_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_30_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_341); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_30_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_344); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_30_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_31_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_352); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_31_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_355); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_31_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_32_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_363); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_32_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_366); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_32_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_33_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_374); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_33_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_377); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_33_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_34_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_385); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_34_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_388); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_34_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_35_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_411); // @[Conditional.scala 40:58 calc6x6.scala 81:22]
  assign Core_35_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_414); // @[Conditional.scala 40:58 calc6x6.scala 82:23]
  assign Core_35_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 80:23]
  assign Core_36_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_283); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_36_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_286); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_36_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_37_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_300); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_37_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_303); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_37_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_38_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_317); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_38_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_320); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_38_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_39_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_331); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_39_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_334); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_39_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_40_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_342); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_40_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_345); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_40_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_41_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_353); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_41_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_356); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_41_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_42_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_364); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_42_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_367); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_42_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_43_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_375); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_43_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_378); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_43_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_44_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_386); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_44_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_389); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_44_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  assign Core_45_io_w_a = _T_2 ? $signed(18'sh0) : $signed(_GEN_412); // @[Conditional.scala 40:58 calc6x6.scala 84:22]
  assign Core_45_io_in_b = _T_2 ? $signed(25'sh0) : $signed(_GEN_415); // @[Conditional.scala 40:58 calc6x6.scala 85:23]
  assign Core_45_io_flag = _T_2 ? 1'h0 : _GEN_278; // @[Conditional.scala 40:58 calc6x6.scala 83:23]
  always @(posedge clock) begin
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_0 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_0 <= {{1{_reg1_mat_real_0_T[16]}},_reg1_mat_real_0_T}; // @[calc6x6.scala 110:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_1 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_1 <= {{1{_reg1_mat_real_1_T[16]}},_reg1_mat_real_1_T}; // @[calc6x6.scala 110:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_2 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_2 <= {{1{_reg1_mat_real_2_T[16]}},_reg1_mat_real_2_T}; // @[calc6x6.scala 110:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_3 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_3 <= {{1{_reg1_mat_real_3_T[16]}},_reg1_mat_real_3_T}; // @[calc6x6.scala 110:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_4 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_4 <= {{1{_reg1_mat_real_4_T[16]}},_reg1_mat_real_4_T}; // @[calc6x6.scala 110:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_5 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_5 <= {{1{_reg1_mat_real_5_T[16]}},_reg1_mat_real_5_T}; // @[calc6x6.scala 110:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_6 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_6 <= _reg1_mat_real_6_T_2[17:0]; // @[calc6x6.scala 111:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_7 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_7 <= _reg1_mat_real_7_T_2[17:0]; // @[calc6x6.scala 111:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_8 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_8 <= _reg1_mat_real_8_T_2[17:0]; // @[calc6x6.scala 111:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_9 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_9 <= _reg1_mat_real_9_T_2[17:0]; // @[calc6x6.scala 111:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_10 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_10 <= _reg1_mat_real_10_T_2[17:0]; // @[calc6x6.scala 111:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_11 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_11 <= _reg1_mat_real_11_T_2[17:0]; // @[calc6x6.scala 111:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_12 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_12 <= _reg1_mat_real_12_T_5[17:0]; // @[calc6x6.scala 112:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_13 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_13 <= _reg1_mat_real_13_T_5[17:0]; // @[calc6x6.scala 112:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_14 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_14 <= _reg1_mat_real_14_T_5[17:0]; // @[calc6x6.scala 112:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_15 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_15 <= _reg1_mat_real_15_T_5[17:0]; // @[calc6x6.scala 112:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_16 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_16 <= _reg1_mat_real_16_T_5[17:0]; // @[calc6x6.scala 112:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_17 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_17 <= _reg1_mat_real_17_T_5[17:0]; // @[calc6x6.scala 112:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_18 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_18 <= {{1{_reg1_mat_real_18_T_3[16]}},_reg1_mat_real_18_T_3}; // @[calc6x6.scala 113:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_19 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_19 <= {{1{_reg1_mat_real_19_T_3[16]}},_reg1_mat_real_19_T_3}; // @[calc6x6.scala 113:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_20 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_20 <= {{1{_reg1_mat_real_20_T_3[16]}},_reg1_mat_real_20_T_3}; // @[calc6x6.scala 113:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_21 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_21 <= {{1{_reg1_mat_real_21_T_3[16]}},_reg1_mat_real_21_T_3}; // @[calc6x6.scala 113:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_22 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_22 <= {{1{_reg1_mat_real_22_T_3[16]}},_reg1_mat_real_22_T_3}; // @[calc6x6.scala 113:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_23 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_23 <= {{1{_reg1_mat_real_23_T_3[16]}},_reg1_mat_real_23_T_3}; // @[calc6x6.scala 113:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_30 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_30 <= {{1{_reg1_mat_real_30_T_3[16]}},_reg1_mat_real_30_T_3}; // @[calc6x6.scala 115:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_31 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_31 <= {{1{_reg1_mat_real_31_T_3[16]}},_reg1_mat_real_31_T_3}; // @[calc6x6.scala 115:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_32 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_32 <= {{1{_reg1_mat_real_32_T_3[16]}},_reg1_mat_real_32_T_3}; // @[calc6x6.scala 115:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_33 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_33 <= {{1{_reg1_mat_real_33_T_3[16]}},_reg1_mat_real_33_T_3}; // @[calc6x6.scala 115:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_34 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_34 <= {{1{_reg1_mat_real_34_T_3[16]}},_reg1_mat_real_34_T_3}; // @[calc6x6.scala 115:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_real_35 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_real_35 <= {{1{_reg1_mat_real_35_T_3[16]}},_reg1_mat_real_35_T_3}; // @[calc6x6.scala 115:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_comp_0 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_comp_0 <= {{1{_reg1_mat_comp_0_T_3[16]}},_reg1_mat_comp_0_T_3}; // @[calc6x6.scala 117:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_comp_1 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_comp_1 <= {{1{_reg1_mat_comp_1_T_3[16]}},_reg1_mat_comp_1_T_3}; // @[calc6x6.scala 117:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_comp_2 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_comp_2 <= {{1{_reg1_mat_comp_2_T_3[16]}},_reg1_mat_comp_2_T_3}; // @[calc6x6.scala 117:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_comp_3 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_comp_3 <= {{1{_reg1_mat_comp_3_T_3[16]}},_reg1_mat_comp_3_T_3}; // @[calc6x6.scala 117:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_comp_4 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_comp_4 <= {{1{_reg1_mat_comp_4_T_3[16]}},_reg1_mat_comp_4_T_3}; // @[calc6x6.scala 117:37]
    end
    if (reset) begin // @[calc6x6.scala 91:23]
      reg1_mat_comp_5 <= 18'sh0; // @[calc6x6.scala 91:23]
    end else begin
      reg1_mat_comp_5 <= {{1{_reg1_mat_comp_5_T_3[16]}},_reg1_mat_comp_5_T_3}; // @[calc6x6.scala 117:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_0 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_0 <= {{1{_reg2_mat_real_0_T[18]}},_reg2_mat_real_0_T}; // @[calc6x6.scala 124:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_1 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_1 <= _reg2_mat_real_1_T_2[19:0]; // @[calc6x6.scala 125:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_2 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_2 <= _reg2_mat_real_2_T_5[19:0]; // @[calc6x6.scala 126:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_3 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_3 <= {{1{_reg2_mat_real_3_T_3[18]}},_reg2_mat_real_3_T_3}; // @[calc6x6.scala 127:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_5 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_5 <= {{1{_reg2_mat_real_5_T_3[18]}},_reg2_mat_real_5_T_3}; // @[calc6x6.scala 129:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_6 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_6 <= {{1{_reg2_mat_real_6_T[18]}},_reg2_mat_real_6_T}; // @[calc6x6.scala 124:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_7 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_7 <= _reg2_mat_real_7_T_2[19:0]; // @[calc6x6.scala 125:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_8 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_8 <= _reg2_mat_real_8_T_5[19:0]; // @[calc6x6.scala 126:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_9 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_9 <= {{1{_reg2_mat_real_9_T_3[18]}},_reg2_mat_real_9_T_3}; // @[calc6x6.scala 127:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_11 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_11 <= {{1{_reg2_mat_real_11_T_3[18]}},_reg2_mat_real_11_T_3}; // @[calc6x6.scala 129:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_12 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_12 <= {{1{_reg2_mat_real_12_T[18]}},_reg2_mat_real_12_T}; // @[calc6x6.scala 124:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_13 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_13 <= _reg2_mat_real_13_T_2[19:0]; // @[calc6x6.scala 125:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_14 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_14 <= _reg2_mat_real_14_T_5[19:0]; // @[calc6x6.scala 126:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_15 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_15 <= {{1{_reg2_mat_real_15_T_3[18]}},_reg2_mat_real_15_T_3}; // @[calc6x6.scala 127:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_17 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_17 <= {{1{_reg2_mat_real_17_T_3[18]}},_reg2_mat_real_17_T_3}; // @[calc6x6.scala 129:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_18 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_18 <= {{1{_reg2_mat_real_18_T[18]}},_reg2_mat_real_18_T}; // @[calc6x6.scala 124:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_19 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_19 <= _reg2_mat_real_19_T_2[19:0]; // @[calc6x6.scala 125:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_20 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_20 <= _reg2_mat_real_20_T_5[19:0]; // @[calc6x6.scala 126:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_21 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_21 <= _reg2_mat_real_21_T_5[19:0]; // @[calc6x6.scala 127:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_22 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_22 <= _reg2_mat_real_22_T_5[19:0]; // @[calc6x6.scala 128:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_23 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_23 <= {{1{_reg2_mat_real_23_T_3[18]}},_reg2_mat_real_23_T_3}; // @[calc6x6.scala 129:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_30 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_30 <= {{1{_reg2_mat_real_30_T[18]}},_reg2_mat_real_30_T}; // @[calc6x6.scala 124:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_31 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_31 <= _reg2_mat_real_31_T_2[19:0]; // @[calc6x6.scala 125:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_32 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_32 <= _reg2_mat_real_32_T_5[19:0]; // @[calc6x6.scala 126:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_33 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_33 <= {{1{_reg2_mat_real_33_T_3[18]}},_reg2_mat_real_33_T_3}; // @[calc6x6.scala 127:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_real_35 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_real_35 <= {{1{_reg2_mat_real_35_T_3[18]}},_reg2_mat_real_35_T_3}; // @[calc6x6.scala 129:37]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_0 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_0 <= {{1{_reg2_mat_comp_0_T[18]}},_reg2_mat_comp_0_T}; // @[calc6x6.scala 132:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_1 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_1 <= _reg2_mat_comp_1_T_2[19:0]; // @[calc6x6.scala 133:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_2 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_2 <= _reg2_mat_comp_2_T_5[19:0]; // @[calc6x6.scala 134:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_3 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_3 <= _reg2_mat_comp_3_T_5[19:0]; // @[calc6x6.scala 135:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_4 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_4 <= _reg2_mat_comp_4_T_5[19:0]; // @[calc6x6.scala 136:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_5 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_5 <= {{1{_reg2_mat_comp_5_T_3[18]}},_reg2_mat_comp_5_T_3}; // @[calc6x6.scala 137:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_6 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_6 <= {{1{_reg2_mat_comp_6_T_3[18]}},_reg2_mat_comp_6_T_3}; // @[calc6x6.scala 140:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_7 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_7 <= {{1{_reg2_mat_comp_7_T_3[18]}},_reg2_mat_comp_7_T_3}; // @[calc6x6.scala 141:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_8 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_8 <= {{1{_reg2_mat_comp_8_T_3[18]}},_reg2_mat_comp_8_T_3}; // @[calc6x6.scala 142:26]
    end
    if (reset) begin // @[calc6x6.scala 92:23]
      reg2_mat_comp_9 <= 20'sh0; // @[calc6x6.scala 92:23]
    end else begin
      reg2_mat_comp_9 <= {{1{_reg2_mat_comp_9_T_3[18]}},_reg2_mat_comp_9_T_3}; // @[calc6x6.scala 143:26]
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_0 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_0 <= _GEN_486[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_1 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_1 <= _GEN_487[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_2 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_2 <= _GEN_488[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_3 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_3 <= _GEN_498[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_4 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_4 <= _GEN_500[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_5 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_5 <= _GEN_502[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_6 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_6 <= _GEN_503[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_7 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_7 <= _GEN_504[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_8 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_8 <= _GEN_505[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_9 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_9 <= _GEN_515[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_10 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_10 <= _GEN_517[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_11 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_11 <= _GEN_519[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_12 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_12 <= _GEN_520[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_13 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_13 <= _GEN_521[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_14 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_14 <= _GEN_522[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_15 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_15 <= _GEN_532[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_16 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_16 <= _GEN_534[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_17 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_17 <= _GEN_536[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_18 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_18 <= _GEN_546[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_19 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_19 <= _GEN_557[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_20 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_20 <= _GEN_568[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_21 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_21 <= _GEN_579[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_22 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_22 <= _GEN_590[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_23 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_23 <= _GEN_601[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_24 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_24 <= _GEN_603[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_25 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_25 <= _GEN_605[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_26 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_26 <= _GEN_607[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_27 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_27 <= _GEN_609[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_28 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_28 <= _GEN_611[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_29 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_29 <= _GEN_613[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_30 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_30 <= _GEN_615[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_31 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_31 <= _GEN_616[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_32 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_32 <= _GEN_617[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_33 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_33 <= _GEN_627[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_34 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_34 <= _GEN_629[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_real_35 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_real_35 <= _GEN_631[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_3 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_3 <= _GEN_499[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_4 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_4 <= _GEN_501[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_9 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_9 <= _GEN_516[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_10 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_10 <= _GEN_518[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_15 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_15 <= _GEN_533[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_16 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_16 <= _GEN_535[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_18 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_18 <= _GEN_547[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_19 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_19 <= _GEN_558[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_20 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_20 <= _GEN_569[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_21 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_21 <= _GEN_580[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_22 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_22 <= _GEN_591[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_23 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_23 <= _GEN_602[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_24 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_24 <= _GEN_604[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_25 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_25 <= _GEN_606[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_26 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_26 <= _GEN_608[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_27 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_27 <= _GEN_610[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_28 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_28 <= _GEN_612[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_29 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_29 <= _GEN_614[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_33 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_33 <= _GEN_628[37:0];
    end
    if (reset) begin // @[calc6x6.scala 93:21]
      w3_mat_comp_34 <= 38'sh0; // @[calc6x6.scala 93:21]
    end else begin
      w3_mat_comp_34 <= _GEN_630[37:0];
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_0 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_0 <= _reg3_mat_real_0_T_12; // @[calc6x6.scala 148:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_1 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_1 <= _reg3_mat_real_1_T_12; // @[calc6x6.scala 148:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_2 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_2 <= _reg3_mat_real_2_T_12; // @[calc6x6.scala 148:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_3 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_3 <= _reg3_mat_real_3_T_12; // @[calc6x6.scala 148:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_4 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_4 <= _reg3_mat_real_4_T_12; // @[calc6x6.scala 148:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_5 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_5 <= _reg3_mat_real_5_T_12; // @[calc6x6.scala 148:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_6 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_6 <= _reg3_mat_real_6_T_9; // @[calc6x6.scala 150:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_7 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_7 <= _reg3_mat_real_7_T_9; // @[calc6x6.scala 150:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_8 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_8 <= _reg3_mat_real_8_T_9; // @[calc6x6.scala 150:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_9 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_9 <= _reg3_mat_real_9_T_9; // @[calc6x6.scala 150:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_10 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_10 <= _reg3_mat_real_10_T_9; // @[calc6x6.scala 150:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_11 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_11 <= _reg3_mat_real_11_T_9; // @[calc6x6.scala 150:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_12 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_12 <= _reg3_mat_real_12_T_9; // @[calc6x6.scala 151:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_13 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_13 <= _reg3_mat_real_13_T_9; // @[calc6x6.scala 151:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_14 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_14 <= _reg3_mat_real_14_T_9; // @[calc6x6.scala 151:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_15 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_15 <= _reg3_mat_real_15_T_9; // @[calc6x6.scala 151:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_16 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_16 <= _reg3_mat_real_16_T_9; // @[calc6x6.scala 151:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_17 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_17 <= _reg3_mat_real_17_T_9; // @[calc6x6.scala 151:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_18 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_18 <= _reg3_mat_real_18_T_12; // @[calc6x6.scala 152:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_19 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_19 <= _reg3_mat_real_19_T_12; // @[calc6x6.scala 152:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_20 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_20 <= _reg3_mat_real_20_T_12; // @[calc6x6.scala 152:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_21 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_21 <= _reg3_mat_real_21_T_12; // @[calc6x6.scala 152:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_22 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_22 <= _reg3_mat_real_22_T_12; // @[calc6x6.scala 152:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_real_23 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_real_23 <= _reg3_mat_real_23_T_12; // @[calc6x6.scala 152:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_comp_3 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_comp_3 <= _reg3_mat_comp_3_T_12; // @[calc6x6.scala 154:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_comp_4 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_comp_4 <= _reg3_mat_comp_4_T_12; // @[calc6x6.scala 154:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_comp_9 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_comp_9 <= _reg3_mat_comp_9_T_9; // @[calc6x6.scala 156:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_comp_10 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_comp_10 <= _reg3_mat_comp_10_T_9; // @[calc6x6.scala 156:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_comp_15 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_comp_15 <= _reg3_mat_comp_15_T_9; // @[calc6x6.scala 157:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_comp_16 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_comp_16 <= _reg3_mat_comp_16_T_9; // @[calc6x6.scala 157:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_comp_21 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_comp_21 <= _reg3_mat_comp_21_T_12; // @[calc6x6.scala 158:37]
    end
    if (reset) begin // @[calc6x6.scala 94:23]
      reg3_mat_comp_22 <= 38'sh0; // @[calc6x6.scala 94:23]
    end else begin
      reg3_mat_comp_22 <= _reg3_mat_comp_22_T_12; // @[calc6x6.scala 158:37]
    end
    if (reset) begin // @[calc6x6.scala 172:28]
      valid_reg_0 <= 1'h0; // @[calc6x6.scala 172:28]
    end else begin
      valid_reg_0 <= io_valid_in; // @[calc6x6.scala 173:18]
    end
    if (reset) begin // @[calc6x6.scala 172:28]
      valid_reg_1 <= 1'h0; // @[calc6x6.scala 172:28]
    end else begin
      valid_reg_1 <= valid_reg_0; // @[calc6x6.scala 175:18]
    end
    if (reset) begin // @[calc6x6.scala 172:28]
      valid_reg_2 <= 1'h0; // @[calc6x6.scala 172:28]
    end else begin
      valid_reg_2 <= valid_reg_1; // @[calc6x6.scala 177:18]
    end
    if (reset) begin // @[calc6x6.scala 172:28]
      valid_reg_3 <= 1'h0; // @[calc6x6.scala 172:28]
    end else begin
      valid_reg_3 <= valid_reg_2; // @[calc6x6.scala 179:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg1_mat_real_0 = _RAND_0[17:0];
  _RAND_1 = {1{`RANDOM}};
  reg1_mat_real_1 = _RAND_1[17:0];
  _RAND_2 = {1{`RANDOM}};
  reg1_mat_real_2 = _RAND_2[17:0];
  _RAND_3 = {1{`RANDOM}};
  reg1_mat_real_3 = _RAND_3[17:0];
  _RAND_4 = {1{`RANDOM}};
  reg1_mat_real_4 = _RAND_4[17:0];
  _RAND_5 = {1{`RANDOM}};
  reg1_mat_real_5 = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  reg1_mat_real_6 = _RAND_6[17:0];
  _RAND_7 = {1{`RANDOM}};
  reg1_mat_real_7 = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  reg1_mat_real_8 = _RAND_8[17:0];
  _RAND_9 = {1{`RANDOM}};
  reg1_mat_real_9 = _RAND_9[17:0];
  _RAND_10 = {1{`RANDOM}};
  reg1_mat_real_10 = _RAND_10[17:0];
  _RAND_11 = {1{`RANDOM}};
  reg1_mat_real_11 = _RAND_11[17:0];
  _RAND_12 = {1{`RANDOM}};
  reg1_mat_real_12 = _RAND_12[17:0];
  _RAND_13 = {1{`RANDOM}};
  reg1_mat_real_13 = _RAND_13[17:0];
  _RAND_14 = {1{`RANDOM}};
  reg1_mat_real_14 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  reg1_mat_real_15 = _RAND_15[17:0];
  _RAND_16 = {1{`RANDOM}};
  reg1_mat_real_16 = _RAND_16[17:0];
  _RAND_17 = {1{`RANDOM}};
  reg1_mat_real_17 = _RAND_17[17:0];
  _RAND_18 = {1{`RANDOM}};
  reg1_mat_real_18 = _RAND_18[17:0];
  _RAND_19 = {1{`RANDOM}};
  reg1_mat_real_19 = _RAND_19[17:0];
  _RAND_20 = {1{`RANDOM}};
  reg1_mat_real_20 = _RAND_20[17:0];
  _RAND_21 = {1{`RANDOM}};
  reg1_mat_real_21 = _RAND_21[17:0];
  _RAND_22 = {1{`RANDOM}};
  reg1_mat_real_22 = _RAND_22[17:0];
  _RAND_23 = {1{`RANDOM}};
  reg1_mat_real_23 = _RAND_23[17:0];
  _RAND_24 = {1{`RANDOM}};
  reg1_mat_real_30 = _RAND_24[17:0];
  _RAND_25 = {1{`RANDOM}};
  reg1_mat_real_31 = _RAND_25[17:0];
  _RAND_26 = {1{`RANDOM}};
  reg1_mat_real_32 = _RAND_26[17:0];
  _RAND_27 = {1{`RANDOM}};
  reg1_mat_real_33 = _RAND_27[17:0];
  _RAND_28 = {1{`RANDOM}};
  reg1_mat_real_34 = _RAND_28[17:0];
  _RAND_29 = {1{`RANDOM}};
  reg1_mat_real_35 = _RAND_29[17:0];
  _RAND_30 = {1{`RANDOM}};
  reg1_mat_comp_0 = _RAND_30[17:0];
  _RAND_31 = {1{`RANDOM}};
  reg1_mat_comp_1 = _RAND_31[17:0];
  _RAND_32 = {1{`RANDOM}};
  reg1_mat_comp_2 = _RAND_32[17:0];
  _RAND_33 = {1{`RANDOM}};
  reg1_mat_comp_3 = _RAND_33[17:0];
  _RAND_34 = {1{`RANDOM}};
  reg1_mat_comp_4 = _RAND_34[17:0];
  _RAND_35 = {1{`RANDOM}};
  reg1_mat_comp_5 = _RAND_35[17:0];
  _RAND_36 = {1{`RANDOM}};
  reg2_mat_real_0 = _RAND_36[19:0];
  _RAND_37 = {1{`RANDOM}};
  reg2_mat_real_1 = _RAND_37[19:0];
  _RAND_38 = {1{`RANDOM}};
  reg2_mat_real_2 = _RAND_38[19:0];
  _RAND_39 = {1{`RANDOM}};
  reg2_mat_real_3 = _RAND_39[19:0];
  _RAND_40 = {1{`RANDOM}};
  reg2_mat_real_5 = _RAND_40[19:0];
  _RAND_41 = {1{`RANDOM}};
  reg2_mat_real_6 = _RAND_41[19:0];
  _RAND_42 = {1{`RANDOM}};
  reg2_mat_real_7 = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  reg2_mat_real_8 = _RAND_43[19:0];
  _RAND_44 = {1{`RANDOM}};
  reg2_mat_real_9 = _RAND_44[19:0];
  _RAND_45 = {1{`RANDOM}};
  reg2_mat_real_11 = _RAND_45[19:0];
  _RAND_46 = {1{`RANDOM}};
  reg2_mat_real_12 = _RAND_46[19:0];
  _RAND_47 = {1{`RANDOM}};
  reg2_mat_real_13 = _RAND_47[19:0];
  _RAND_48 = {1{`RANDOM}};
  reg2_mat_real_14 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  reg2_mat_real_15 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  reg2_mat_real_17 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  reg2_mat_real_18 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  reg2_mat_real_19 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  reg2_mat_real_20 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  reg2_mat_real_21 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  reg2_mat_real_22 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  reg2_mat_real_23 = _RAND_56[19:0];
  _RAND_57 = {1{`RANDOM}};
  reg2_mat_real_30 = _RAND_57[19:0];
  _RAND_58 = {1{`RANDOM}};
  reg2_mat_real_31 = _RAND_58[19:0];
  _RAND_59 = {1{`RANDOM}};
  reg2_mat_real_32 = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  reg2_mat_real_33 = _RAND_60[19:0];
  _RAND_61 = {1{`RANDOM}};
  reg2_mat_real_35 = _RAND_61[19:0];
  _RAND_62 = {1{`RANDOM}};
  reg2_mat_comp_0 = _RAND_62[19:0];
  _RAND_63 = {1{`RANDOM}};
  reg2_mat_comp_1 = _RAND_63[19:0];
  _RAND_64 = {1{`RANDOM}};
  reg2_mat_comp_2 = _RAND_64[19:0];
  _RAND_65 = {1{`RANDOM}};
  reg2_mat_comp_3 = _RAND_65[19:0];
  _RAND_66 = {1{`RANDOM}};
  reg2_mat_comp_4 = _RAND_66[19:0];
  _RAND_67 = {1{`RANDOM}};
  reg2_mat_comp_5 = _RAND_67[19:0];
  _RAND_68 = {1{`RANDOM}};
  reg2_mat_comp_6 = _RAND_68[19:0];
  _RAND_69 = {1{`RANDOM}};
  reg2_mat_comp_7 = _RAND_69[19:0];
  _RAND_70 = {1{`RANDOM}};
  reg2_mat_comp_8 = _RAND_70[19:0];
  _RAND_71 = {1{`RANDOM}};
  reg2_mat_comp_9 = _RAND_71[19:0];
  _RAND_72 = {2{`RANDOM}};
  w3_mat_real_0 = _RAND_72[37:0];
  _RAND_73 = {2{`RANDOM}};
  w3_mat_real_1 = _RAND_73[37:0];
  _RAND_74 = {2{`RANDOM}};
  w3_mat_real_2 = _RAND_74[37:0];
  _RAND_75 = {2{`RANDOM}};
  w3_mat_real_3 = _RAND_75[37:0];
  _RAND_76 = {2{`RANDOM}};
  w3_mat_real_4 = _RAND_76[37:0];
  _RAND_77 = {2{`RANDOM}};
  w3_mat_real_5 = _RAND_77[37:0];
  _RAND_78 = {2{`RANDOM}};
  w3_mat_real_6 = _RAND_78[37:0];
  _RAND_79 = {2{`RANDOM}};
  w3_mat_real_7 = _RAND_79[37:0];
  _RAND_80 = {2{`RANDOM}};
  w3_mat_real_8 = _RAND_80[37:0];
  _RAND_81 = {2{`RANDOM}};
  w3_mat_real_9 = _RAND_81[37:0];
  _RAND_82 = {2{`RANDOM}};
  w3_mat_real_10 = _RAND_82[37:0];
  _RAND_83 = {2{`RANDOM}};
  w3_mat_real_11 = _RAND_83[37:0];
  _RAND_84 = {2{`RANDOM}};
  w3_mat_real_12 = _RAND_84[37:0];
  _RAND_85 = {2{`RANDOM}};
  w3_mat_real_13 = _RAND_85[37:0];
  _RAND_86 = {2{`RANDOM}};
  w3_mat_real_14 = _RAND_86[37:0];
  _RAND_87 = {2{`RANDOM}};
  w3_mat_real_15 = _RAND_87[37:0];
  _RAND_88 = {2{`RANDOM}};
  w3_mat_real_16 = _RAND_88[37:0];
  _RAND_89 = {2{`RANDOM}};
  w3_mat_real_17 = _RAND_89[37:0];
  _RAND_90 = {2{`RANDOM}};
  w3_mat_real_18 = _RAND_90[37:0];
  _RAND_91 = {2{`RANDOM}};
  w3_mat_real_19 = _RAND_91[37:0];
  _RAND_92 = {2{`RANDOM}};
  w3_mat_real_20 = _RAND_92[37:0];
  _RAND_93 = {2{`RANDOM}};
  w3_mat_real_21 = _RAND_93[37:0];
  _RAND_94 = {2{`RANDOM}};
  w3_mat_real_22 = _RAND_94[37:0];
  _RAND_95 = {2{`RANDOM}};
  w3_mat_real_23 = _RAND_95[37:0];
  _RAND_96 = {2{`RANDOM}};
  w3_mat_real_24 = _RAND_96[37:0];
  _RAND_97 = {2{`RANDOM}};
  w3_mat_real_25 = _RAND_97[37:0];
  _RAND_98 = {2{`RANDOM}};
  w3_mat_real_26 = _RAND_98[37:0];
  _RAND_99 = {2{`RANDOM}};
  w3_mat_real_27 = _RAND_99[37:0];
  _RAND_100 = {2{`RANDOM}};
  w3_mat_real_28 = _RAND_100[37:0];
  _RAND_101 = {2{`RANDOM}};
  w3_mat_real_29 = _RAND_101[37:0];
  _RAND_102 = {2{`RANDOM}};
  w3_mat_real_30 = _RAND_102[37:0];
  _RAND_103 = {2{`RANDOM}};
  w3_mat_real_31 = _RAND_103[37:0];
  _RAND_104 = {2{`RANDOM}};
  w3_mat_real_32 = _RAND_104[37:0];
  _RAND_105 = {2{`RANDOM}};
  w3_mat_real_33 = _RAND_105[37:0];
  _RAND_106 = {2{`RANDOM}};
  w3_mat_real_34 = _RAND_106[37:0];
  _RAND_107 = {2{`RANDOM}};
  w3_mat_real_35 = _RAND_107[37:0];
  _RAND_108 = {2{`RANDOM}};
  w3_mat_comp_3 = _RAND_108[37:0];
  _RAND_109 = {2{`RANDOM}};
  w3_mat_comp_4 = _RAND_109[37:0];
  _RAND_110 = {2{`RANDOM}};
  w3_mat_comp_9 = _RAND_110[37:0];
  _RAND_111 = {2{`RANDOM}};
  w3_mat_comp_10 = _RAND_111[37:0];
  _RAND_112 = {2{`RANDOM}};
  w3_mat_comp_15 = _RAND_112[37:0];
  _RAND_113 = {2{`RANDOM}};
  w3_mat_comp_16 = _RAND_113[37:0];
  _RAND_114 = {2{`RANDOM}};
  w3_mat_comp_18 = _RAND_114[37:0];
  _RAND_115 = {2{`RANDOM}};
  w3_mat_comp_19 = _RAND_115[37:0];
  _RAND_116 = {2{`RANDOM}};
  w3_mat_comp_20 = _RAND_116[37:0];
  _RAND_117 = {2{`RANDOM}};
  w3_mat_comp_21 = _RAND_117[37:0];
  _RAND_118 = {2{`RANDOM}};
  w3_mat_comp_22 = _RAND_118[37:0];
  _RAND_119 = {2{`RANDOM}};
  w3_mat_comp_23 = _RAND_119[37:0];
  _RAND_120 = {2{`RANDOM}};
  w3_mat_comp_24 = _RAND_120[37:0];
  _RAND_121 = {2{`RANDOM}};
  w3_mat_comp_25 = _RAND_121[37:0];
  _RAND_122 = {2{`RANDOM}};
  w3_mat_comp_26 = _RAND_122[37:0];
  _RAND_123 = {2{`RANDOM}};
  w3_mat_comp_27 = _RAND_123[37:0];
  _RAND_124 = {2{`RANDOM}};
  w3_mat_comp_28 = _RAND_124[37:0];
  _RAND_125 = {2{`RANDOM}};
  w3_mat_comp_29 = _RAND_125[37:0];
  _RAND_126 = {2{`RANDOM}};
  w3_mat_comp_33 = _RAND_126[37:0];
  _RAND_127 = {2{`RANDOM}};
  w3_mat_comp_34 = _RAND_127[37:0];
  _RAND_128 = {2{`RANDOM}};
  reg3_mat_real_0 = _RAND_128[37:0];
  _RAND_129 = {2{`RANDOM}};
  reg3_mat_real_1 = _RAND_129[37:0];
  _RAND_130 = {2{`RANDOM}};
  reg3_mat_real_2 = _RAND_130[37:0];
  _RAND_131 = {2{`RANDOM}};
  reg3_mat_real_3 = _RAND_131[37:0];
  _RAND_132 = {2{`RANDOM}};
  reg3_mat_real_4 = _RAND_132[37:0];
  _RAND_133 = {2{`RANDOM}};
  reg3_mat_real_5 = _RAND_133[37:0];
  _RAND_134 = {2{`RANDOM}};
  reg3_mat_real_6 = _RAND_134[37:0];
  _RAND_135 = {2{`RANDOM}};
  reg3_mat_real_7 = _RAND_135[37:0];
  _RAND_136 = {2{`RANDOM}};
  reg3_mat_real_8 = _RAND_136[37:0];
  _RAND_137 = {2{`RANDOM}};
  reg3_mat_real_9 = _RAND_137[37:0];
  _RAND_138 = {2{`RANDOM}};
  reg3_mat_real_10 = _RAND_138[37:0];
  _RAND_139 = {2{`RANDOM}};
  reg3_mat_real_11 = _RAND_139[37:0];
  _RAND_140 = {2{`RANDOM}};
  reg3_mat_real_12 = _RAND_140[37:0];
  _RAND_141 = {2{`RANDOM}};
  reg3_mat_real_13 = _RAND_141[37:0];
  _RAND_142 = {2{`RANDOM}};
  reg3_mat_real_14 = _RAND_142[37:0];
  _RAND_143 = {2{`RANDOM}};
  reg3_mat_real_15 = _RAND_143[37:0];
  _RAND_144 = {2{`RANDOM}};
  reg3_mat_real_16 = _RAND_144[37:0];
  _RAND_145 = {2{`RANDOM}};
  reg3_mat_real_17 = _RAND_145[37:0];
  _RAND_146 = {2{`RANDOM}};
  reg3_mat_real_18 = _RAND_146[37:0];
  _RAND_147 = {2{`RANDOM}};
  reg3_mat_real_19 = _RAND_147[37:0];
  _RAND_148 = {2{`RANDOM}};
  reg3_mat_real_20 = _RAND_148[37:0];
  _RAND_149 = {2{`RANDOM}};
  reg3_mat_real_21 = _RAND_149[37:0];
  _RAND_150 = {2{`RANDOM}};
  reg3_mat_real_22 = _RAND_150[37:0];
  _RAND_151 = {2{`RANDOM}};
  reg3_mat_real_23 = _RAND_151[37:0];
  _RAND_152 = {2{`RANDOM}};
  reg3_mat_comp_3 = _RAND_152[37:0];
  _RAND_153 = {2{`RANDOM}};
  reg3_mat_comp_4 = _RAND_153[37:0];
  _RAND_154 = {2{`RANDOM}};
  reg3_mat_comp_9 = _RAND_154[37:0];
  _RAND_155 = {2{`RANDOM}};
  reg3_mat_comp_10 = _RAND_155[37:0];
  _RAND_156 = {2{`RANDOM}};
  reg3_mat_comp_15 = _RAND_156[37:0];
  _RAND_157 = {2{`RANDOM}};
  reg3_mat_comp_16 = _RAND_157[37:0];
  _RAND_158 = {2{`RANDOM}};
  reg3_mat_comp_21 = _RAND_158[37:0];
  _RAND_159 = {2{`RANDOM}};
  reg3_mat_comp_22 = _RAND_159[37:0];
  _RAND_160 = {1{`RANDOM}};
  valid_reg_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_reg_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_reg_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_reg_3 = _RAND_163[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Calc8x8(
  input         clock,
  input         reset,
  input  [15:0] io_input_mat_0,
  input  [15:0] io_input_mat_1,
  input  [15:0] io_input_mat_2,
  input  [15:0] io_input_mat_3,
  input  [15:0] io_input_mat_4,
  input  [15:0] io_input_mat_5,
  input  [15:0] io_input_mat_6,
  input  [15:0] io_input_mat_7,
  input  [15:0] io_input_mat_8,
  input  [15:0] io_input_mat_9,
  input  [15:0] io_input_mat_10,
  input  [15:0] io_input_mat_11,
  input  [15:0] io_input_mat_12,
  input  [15:0] io_input_mat_13,
  input  [15:0] io_input_mat_14,
  input  [15:0] io_input_mat_15,
  input  [15:0] io_input_mat_16,
  input  [15:0] io_input_mat_17,
  input  [15:0] io_input_mat_18,
  input  [15:0] io_input_mat_19,
  input  [15:0] io_input_mat_20,
  input  [15:0] io_input_mat_21,
  input  [15:0] io_input_mat_22,
  input  [15:0] io_input_mat_23,
  input  [15:0] io_input_mat_24,
  input  [15:0] io_input_mat_25,
  input  [15:0] io_input_mat_26,
  input  [15:0] io_input_mat_27,
  input  [15:0] io_input_mat_28,
  input  [15:0] io_input_mat_29,
  input  [15:0] io_input_mat_30,
  input  [15:0] io_input_mat_31,
  input  [15:0] io_input_mat_32,
  input  [15:0] io_input_mat_33,
  input  [15:0] io_input_mat_34,
  input  [15:0] io_input_mat_35,
  input  [15:0] io_input_mat_36,
  input  [15:0] io_input_mat_37,
  input  [15:0] io_input_mat_38,
  input  [15:0] io_input_mat_39,
  input  [15:0] io_input_mat_40,
  input  [15:0] io_input_mat_41,
  input  [15:0] io_input_mat_42,
  input  [15:0] io_input_mat_43,
  input  [15:0] io_input_mat_44,
  input  [15:0] io_input_mat_45,
  input  [15:0] io_input_mat_46,
  input  [15:0] io_input_mat_47,
  input  [15:0] io_input_mat_48,
  input  [15:0] io_input_mat_49,
  input  [15:0] io_input_mat_50,
  input  [15:0] io_input_mat_51,
  input  [15:0] io_input_mat_52,
  input  [15:0] io_input_mat_53,
  input  [15:0] io_input_mat_54,
  input  [15:0] io_input_mat_55,
  input  [15:0] io_input_mat_56,
  input  [15:0] io_input_mat_57,
  input  [15:0] io_input_mat_58,
  input  [15:0] io_input_mat_59,
  input  [15:0] io_input_mat_60,
  input  [15:0] io_input_mat_61,
  input  [15:0] io_input_mat_62,
  input  [15:0] io_input_mat_63,
  input  [15:0] io_input_up_0,
  input  [15:0] io_input_up_1,
  input  [15:0] io_input_up_2,
  input  [15:0] io_input_up_3,
  input  [15:0] io_input_up_4,
  input  [15:0] io_input_up_5,
  input  [15:0] io_input_up_6,
  input  [15:0] io_input_up_7,
  input  [15:0] io_input_up_8,
  input  [15:0] io_input_up_9,
  input  [15:0] io_input_down_0,
  input  [15:0] io_input_down_1,
  input  [15:0] io_input_down_2,
  input  [15:0] io_input_down_3,
  input  [15:0] io_input_down_4,
  input  [15:0] io_input_down_5,
  input  [15:0] io_input_down_6,
  input  [15:0] io_input_down_7,
  input  [15:0] io_input_down_8,
  input  [15:0] io_input_down_9,
  input  [15:0] io_input_left_0,
  input  [15:0] io_input_left_1,
  input  [15:0] io_input_left_2,
  input  [15:0] io_input_left_3,
  input  [15:0] io_input_left_4,
  input  [15:0] io_input_left_5,
  input  [15:0] io_input_left_6,
  input  [15:0] io_input_left_7,
  input  [15:0] io_input_right_0,
  input  [15:0] io_input_right_1,
  input  [15:0] io_input_right_2,
  input  [15:0] io_input_right_3,
  input  [15:0] io_input_right_4,
  input  [15:0] io_input_right_5,
  input  [15:0] io_input_right_6,
  input  [15:0] io_input_right_7,
  input  [1:0]  io_flag,
  input  [15:0] io_weight_0_real_0,
  input  [15:0] io_weight_0_real_1,
  input  [15:0] io_weight_0_real_2,
  input  [15:0] io_weight_0_real_3,
  input  [15:0] io_weight_0_real_4,
  input  [15:0] io_weight_0_real_5,
  input  [15:0] io_weight_0_real_6,
  input  [15:0] io_weight_0_real_7,
  input  [15:0] io_weight_0_real_8,
  input  [15:0] io_weight_0_real_9,
  input  [15:0] io_weight_0_real_10,
  input  [15:0] io_weight_0_real_11,
  input  [15:0] io_weight_0_real_12,
  input  [15:0] io_weight_0_real_13,
  input  [15:0] io_weight_0_real_14,
  input  [15:0] io_weight_0_real_15,
  input  [15:0] io_weight_1_real_0,
  input  [15:0] io_weight_1_real_1,
  input  [15:0] io_weight_1_real_2,
  input  [15:0] io_weight_1_real_3,
  input  [15:0] io_weight_1_real_4,
  input  [15:0] io_weight_1_real_5,
  input  [15:0] io_weight_1_real_6,
  input  [15:0] io_weight_1_real_7,
  input  [15:0] io_weight_1_real_8,
  input  [15:0] io_weight_1_real_9,
  input  [15:0] io_weight_1_real_10,
  input  [15:0] io_weight_1_real_11,
  input  [15:0] io_weight_1_real_12,
  input  [15:0] io_weight_1_real_13,
  input  [15:0] io_weight_1_real_14,
  input  [15:0] io_weight_1_real_15,
  input  [15:0] io_weight_2_real_0,
  input  [15:0] io_weight_2_real_1,
  input  [15:0] io_weight_2_real_2,
  input  [15:0] io_weight_2_real_3,
  input  [15:0] io_weight_2_real_4,
  input  [15:0] io_weight_2_real_5,
  input  [15:0] io_weight_2_real_6,
  input  [15:0] io_weight_2_real_7,
  input  [15:0] io_weight_2_real_8,
  input  [15:0] io_weight_2_real_9,
  input  [15:0] io_weight_2_real_10,
  input  [15:0] io_weight_2_real_11,
  input  [15:0] io_weight_2_real_12,
  input  [15:0] io_weight_2_real_13,
  input  [15:0] io_weight_2_real_14,
  input  [15:0] io_weight_2_real_15,
  input  [15:0] io_weight_3_real_0,
  input  [15:0] io_weight_3_real_1,
  input  [15:0] io_weight_3_real_2,
  input  [15:0] io_weight_3_real_3,
  input  [15:0] io_weight_3_real_4,
  input  [15:0] io_weight_3_real_5,
  input  [15:0] io_weight_3_real_6,
  input  [15:0] io_weight_3_real_7,
  input  [15:0] io_weight_3_real_8,
  input  [15:0] io_weight_3_real_9,
  input  [15:0] io_weight_3_real_10,
  input  [15:0] io_weight_3_real_11,
  input  [15:0] io_weight_3_real_12,
  input  [15:0] io_weight_3_real_13,
  input  [15:0] io_weight_3_real_14,
  input  [15:0] io_weight_3_real_15,
  output [36:0] io_output_mat_0,
  output [36:0] io_output_mat_1,
  output [36:0] io_output_mat_2,
  output [36:0] io_output_mat_3,
  output [36:0] io_output_mat_4,
  output [36:0] io_output_mat_5,
  output [36:0] io_output_mat_6,
  output [36:0] io_output_mat_7,
  output [36:0] io_output_mat_8,
  output [36:0] io_output_mat_9,
  output [36:0] io_output_mat_10,
  output [36:0] io_output_mat_11,
  output [36:0] io_output_mat_12,
  output [36:0] io_output_mat_13,
  output [36:0] io_output_mat_14,
  output [36:0] io_output_mat_15,
  output [36:0] io_output_mat_16,
  output [36:0] io_output_mat_17,
  output [36:0] io_output_mat_18,
  output [36:0] io_output_mat_19,
  output [36:0] io_output_mat_20,
  output [36:0] io_output_mat_21,
  output [36:0] io_output_mat_22,
  output [36:0] io_output_mat_23,
  output [36:0] io_output_mat_24,
  output [36:0] io_output_mat_25,
  output [36:0] io_output_mat_26,
  output [36:0] io_output_mat_27,
  output [36:0] io_output_mat_28,
  output [36:0] io_output_mat_29,
  output [36:0] io_output_mat_30,
  output [36:0] io_output_mat_31,
  output [36:0] io_output_mat_32,
  output [36:0] io_output_mat_33,
  output [36:0] io_output_mat_34,
  output [36:0] io_output_mat_35,
  output [36:0] io_output_mat_36,
  output [36:0] io_output_mat_37,
  output [36:0] io_output_mat_38,
  output [36:0] io_output_mat_39,
  output [36:0] io_output_mat_40,
  output [36:0] io_output_mat_41,
  output [36:0] io_output_mat_42,
  output [36:0] io_output_mat_43,
  output [36:0] io_output_mat_44,
  output [36:0] io_output_mat_45,
  output [36:0] io_output_mat_46,
  output [36:0] io_output_mat_47,
  output [36:0] io_output_mat_48,
  output [36:0] io_output_mat_49,
  output [36:0] io_output_mat_50,
  output [36:0] io_output_mat_51,
  output [36:0] io_output_mat_52,
  output [36:0] io_output_mat_53,
  output [36:0] io_output_mat_54,
  output [36:0] io_output_mat_55,
  output [36:0] io_output_mat_56,
  output [36:0] io_output_mat_57,
  output [36:0] io_output_mat_58,
  output [36:0] io_output_mat_59,
  output [36:0] io_output_mat_60,
  output [36:0] io_output_mat_61,
  output [36:0] io_output_mat_62,
  output [36:0] io_output_mat_63,
  input         io_valid_in,
  output        io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
`endif // RANDOMIZE_REG_INIT
  wire  Calc6x6_clock; // @[calc8x8.scala 59:39]
  wire  Calc6x6_reset; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_0; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_1; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_2; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_3; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_4; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_5; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_6; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_7; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_8; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_9; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_10; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_11; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_12; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_13; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_14; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_15; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_16; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_17; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_18; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_19; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_20; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_21; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_22; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_23; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_24; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_25; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_26; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_27; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_28; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_29; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_30; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_31; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_32; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_33; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_34; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_io_input_mat_35; // @[calc8x8.scala 59:39]
  wire [1:0] Calc6x6_io_flag; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_10; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_11; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_12; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_13; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_14; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_real_15; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp1_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp2_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_io_weight_comp3_9; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_0; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_1; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_2; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_3; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_4; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_5; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_6; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_7; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_8; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_9; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_10; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_11; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_12; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_13; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_14; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_io_output_mat_15; // @[calc8x8.scala 59:39]
  wire  Calc6x6_io_valid_in; // @[calc8x8.scala 59:39]
  wire  Calc6x6_io_valid_out; // @[calc8x8.scala 59:39]
  wire  Calc6x6_1_clock; // @[calc8x8.scala 59:39]
  wire  Calc6x6_1_reset; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_0; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_1; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_2; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_3; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_4; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_5; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_6; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_7; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_8; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_9; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_10; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_11; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_12; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_13; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_14; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_15; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_16; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_17; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_18; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_19; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_20; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_21; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_22; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_23; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_24; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_25; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_26; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_27; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_28; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_29; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_30; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_31; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_32; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_33; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_34; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_1_io_input_mat_35; // @[calc8x8.scala 59:39]
  wire [1:0] Calc6x6_1_io_flag; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_10; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_11; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_12; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_13; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_14; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_real_15; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp1_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp2_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_1_io_weight_comp3_9; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_0; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_1; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_2; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_3; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_4; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_5; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_6; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_7; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_8; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_9; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_10; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_11; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_12; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_13; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_14; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_1_io_output_mat_15; // @[calc8x8.scala 59:39]
  wire  Calc6x6_1_io_valid_in; // @[calc8x8.scala 59:39]
  wire  Calc6x6_1_io_valid_out; // @[calc8x8.scala 59:39]
  wire  Calc6x6_2_clock; // @[calc8x8.scala 59:39]
  wire  Calc6x6_2_reset; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_0; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_1; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_2; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_3; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_4; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_5; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_6; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_7; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_8; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_9; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_10; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_11; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_12; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_13; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_14; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_15; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_16; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_17; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_18; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_19; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_20; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_21; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_22; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_23; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_24; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_25; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_26; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_27; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_28; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_29; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_30; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_31; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_32; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_33; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_34; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_2_io_input_mat_35; // @[calc8x8.scala 59:39]
  wire [1:0] Calc6x6_2_io_flag; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_10; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_11; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_12; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_13; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_14; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_real_15; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp1_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp2_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_2_io_weight_comp3_9; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_0; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_1; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_2; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_3; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_4; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_5; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_6; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_7; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_8; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_9; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_10; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_11; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_12; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_13; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_14; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_2_io_output_mat_15; // @[calc8x8.scala 59:39]
  wire  Calc6x6_2_io_valid_in; // @[calc8x8.scala 59:39]
  wire  Calc6x6_2_io_valid_out; // @[calc8x8.scala 59:39]
  wire  Calc6x6_3_clock; // @[calc8x8.scala 59:39]
  wire  Calc6x6_3_reset; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_0; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_1; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_2; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_3; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_4; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_5; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_6; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_7; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_8; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_9; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_10; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_11; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_12; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_13; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_14; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_15; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_16; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_17; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_18; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_19; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_20; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_21; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_22; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_23; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_24; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_25; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_26; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_27; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_28; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_29; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_30; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_31; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_32; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_33; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_34; // @[calc8x8.scala 59:39]
  wire [15:0] Calc6x6_3_io_input_mat_35; // @[calc8x8.scala 59:39]
  wire [1:0] Calc6x6_3_io_flag; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_10; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_11; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_12; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_13; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_14; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_real_15; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp1_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp2_9; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_0; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_1; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_2; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_3; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_4; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_5; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_6; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_7; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_8; // @[calc8x8.scala 59:39]
  wire [17:0] Calc6x6_3_io_weight_comp3_9; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_0; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_1; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_2; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_3; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_4; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_5; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_6; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_7; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_8; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_9; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_10; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_11; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_12; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_13; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_14; // @[calc8x8.scala 59:39]
  wire [36:0] Calc6x6_3_io_output_mat_15; // @[calc8x8.scala 59:39]
  wire  Calc6x6_3_io_valid_in; // @[calc8x8.scala 59:39]
  wire  Calc6x6_3_io_valid_out; // @[calc8x8.scala 59:39]
  reg [17:0] _B_0_0; // @[calc8x8.scala 71:21]
  reg [17:0] _B_0_1; // @[calc8x8.scala 71:21]
  reg [17:0] _B_0_2; // @[calc8x8.scala 71:21]
  reg [17:0] _B_1_0; // @[calc8x8.scala 71:21]
  reg [17:0] _B_1_1; // @[calc8x8.scala 71:21]
  reg [17:0] _B_1_2; // @[calc8x8.scala 71:21]
  reg [17:0] _B_2_0; // @[calc8x8.scala 71:21]
  reg [17:0] _B_2_1; // @[calc8x8.scala 71:21]
  reg [17:0] _B_2_2; // @[calc8x8.scala 71:21]
  reg [17:0] _B_3_0; // @[calc8x8.scala 71:21]
  reg [17:0] _B_3_1; // @[calc8x8.scala 71:21]
  reg [17:0] _B_3_2; // @[calc8x8.scala 71:21]
  reg [17:0] _B_5_0; // @[calc8x8.scala 71:21]
  reg [17:0] _B_5_1; // @[calc8x8.scala 71:21]
  reg [17:0] _B_5_2; // @[calc8x8.scala 71:21]
  reg [17:0] _Bi_3_0; // @[calc8x8.scala 72:22]
  reg [17:0] _Bi_3_1; // @[calc8x8.scala 72:22]
  reg [17:0] _Bi_3_2; // @[calc8x8.scala 72:22]
  wire [15:0] __B_1_0_T_2 = $signed(io_weight_0_real_0) + $signed(io_weight_0_real_3); // @[calc8x8.scala 79:28]
  wire [15:0] __B_1_0_T_5 = $signed(__B_1_0_T_2) + $signed(io_weight_0_real_6); // @[calc8x8.scala 79:36]
  wire [15:0] __B_2_0_T_2 = $signed(io_weight_0_real_0) - $signed(io_weight_0_real_3); // @[calc8x8.scala 80:28]
  wire [15:0] __B_2_0_T_5 = $signed(__B_2_0_T_2) + $signed(io_weight_0_real_6); // @[calc8x8.scala 80:36]
  wire [15:0] __B_3_0_T_2 = $signed(io_weight_0_real_0) - $signed(io_weight_0_real_6); // @[calc8x8.scala 81:28]
  wire [15:0] __B_1_1_T_2 = $signed(io_weight_0_real_1) + $signed(io_weight_0_real_4); // @[calc8x8.scala 79:28]
  wire [15:0] __B_1_1_T_5 = $signed(__B_1_1_T_2) + $signed(io_weight_0_real_7); // @[calc8x8.scala 79:36]
  wire [15:0] __B_2_1_T_2 = $signed(io_weight_0_real_1) - $signed(io_weight_0_real_4); // @[calc8x8.scala 80:28]
  wire [15:0] __B_2_1_T_5 = $signed(__B_2_1_T_2) + $signed(io_weight_0_real_7); // @[calc8x8.scala 80:36]
  wire [15:0] __B_3_1_T_2 = $signed(io_weight_0_real_1) - $signed(io_weight_0_real_7); // @[calc8x8.scala 81:28]
  wire [15:0] __B_1_2_T_2 = $signed(io_weight_0_real_2) + $signed(io_weight_0_real_5); // @[calc8x8.scala 79:28]
  wire [15:0] __B_1_2_T_5 = $signed(__B_1_2_T_2) + $signed(io_weight_0_real_8); // @[calc8x8.scala 79:36]
  wire [15:0] __B_2_2_T_2 = $signed(io_weight_0_real_2) - $signed(io_weight_0_real_5); // @[calc8x8.scala 80:28]
  wire [15:0] __B_2_2_T_5 = $signed(__B_2_2_T_2) + $signed(io_weight_0_real_8); // @[calc8x8.scala 80:36]
  wire [15:0] __B_3_2_T_2 = $signed(io_weight_0_real_2) - $signed(io_weight_0_real_8); // @[calc8x8.scala 81:28]
  reg [18:0] __B_0_0; // @[calc8x8.scala 89:22]
  reg [18:0] __B_0_1; // @[calc8x8.scala 89:22]
  reg [18:0] __B_0_2; // @[calc8x8.scala 89:22]
  reg [18:0] __B_0_3; // @[calc8x8.scala 89:22]
  reg [18:0] __B_0_5; // @[calc8x8.scala 89:22]
  reg [18:0] __B_1_0; // @[calc8x8.scala 89:22]
  reg [18:0] __B_1_1; // @[calc8x8.scala 89:22]
  reg [18:0] __B_1_2; // @[calc8x8.scala 89:22]
  reg [18:0] __B_1_3; // @[calc8x8.scala 89:22]
  reg [18:0] __B_1_5; // @[calc8x8.scala 89:22]
  reg [18:0] __B_2_0; // @[calc8x8.scala 89:22]
  reg [18:0] __B_2_1; // @[calc8x8.scala 89:22]
  reg [18:0] __B_2_2; // @[calc8x8.scala 89:22]
  reg [18:0] __B_2_3; // @[calc8x8.scala 89:22]
  reg [18:0] __B_2_5; // @[calc8x8.scala 89:22]
  reg [18:0] __B_3_0; // @[calc8x8.scala 89:22]
  reg [18:0] __B_3_1; // @[calc8x8.scala 89:22]
  reg [18:0] __B_3_2; // @[calc8x8.scala 89:22]
  reg [18:0] __B_3_3; // @[calc8x8.scala 89:22]
  reg [18:0] __B_3_4; // @[calc8x8.scala 89:22]
  reg [18:0] __B_3_5; // @[calc8x8.scala 89:22]
  reg [18:0] __B_5_0; // @[calc8x8.scala 89:22]
  reg [18:0] __B_5_1; // @[calc8x8.scala 89:22]
  reg [18:0] __B_5_2; // @[calc8x8.scala 89:22]
  reg [18:0] __B_5_3; // @[calc8x8.scala 89:22]
  reg [18:0] __B_5_5; // @[calc8x8.scala 89:22]
  reg [18:0] __Bi_0_3; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_1_3; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_2_3; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_3_0; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_3_1; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_3_2; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_3_3; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_3_4; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_3_5; // @[calc8x8.scala 90:23]
  reg [18:0] __Bi_5_3; // @[calc8x8.scala 90:23]
  wire [17:0] ___B_0_1_T_2 = $signed(_B_0_0) + $signed(_B_0_1); // @[calc8x8.scala 94:30]
  wire [17:0] ___B_0_1_T_5 = $signed(___B_0_1_T_2) + $signed(_B_0_2); // @[calc8x8.scala 94:39]
  wire [17:0] ___B_0_2_T_2 = $signed(_B_0_0) - $signed(_B_0_1); // @[calc8x8.scala 95:30]
  wire [17:0] ___B_0_2_T_5 = $signed(___B_0_2_T_2) + $signed(_B_0_2); // @[calc8x8.scala 95:39]
  wire [17:0] ___B_0_3_T_2 = $signed(_B_0_0) - $signed(_B_0_2); // @[calc8x8.scala 96:30]
  wire [17:0] ___B_0_3_T_5 = $signed(___B_0_3_T_2) - 18'sh0; // @[calc8x8.scala 96:39]
  wire [18:0] ___Bi_0_3_T_3 = {{1{_B_0_1[17]}},_B_0_1}; // @[calc8x8.scala 102:42]
  wire [17:0] ___Bi_0_3_T_5 = ___Bi_0_3_T_3[17:0]; // @[calc8x8.scala 102:42]
  wire [17:0] ___B_1_1_T_2 = $signed(_B_1_0) + $signed(_B_1_1); // @[calc8x8.scala 94:30]
  wire [17:0] ___B_1_1_T_5 = $signed(___B_1_1_T_2) + $signed(_B_1_2); // @[calc8x8.scala 94:39]
  wire [17:0] ___B_1_2_T_2 = $signed(_B_1_0) - $signed(_B_1_1); // @[calc8x8.scala 95:30]
  wire [17:0] ___B_1_2_T_5 = $signed(___B_1_2_T_2) + $signed(_B_1_2); // @[calc8x8.scala 95:39]
  wire [17:0] ___B_1_3_T_2 = $signed(_B_1_0) - $signed(_B_1_2); // @[calc8x8.scala 96:30]
  wire [17:0] ___B_1_3_T_5 = $signed(___B_1_3_T_2) - 18'sh0; // @[calc8x8.scala 96:39]
  wire [18:0] ___Bi_1_3_T_3 = {{1{_B_1_1[17]}},_B_1_1}; // @[calc8x8.scala 102:42]
  wire [17:0] ___Bi_1_3_T_5 = ___Bi_1_3_T_3[17:0]; // @[calc8x8.scala 102:42]
  wire [17:0] ___B_2_1_T_2 = $signed(_B_2_0) + $signed(_B_2_1); // @[calc8x8.scala 94:30]
  wire [17:0] ___B_2_1_T_5 = $signed(___B_2_1_T_2) + $signed(_B_2_2); // @[calc8x8.scala 94:39]
  wire [17:0] ___B_2_2_T_2 = $signed(_B_2_0) - $signed(_B_2_1); // @[calc8x8.scala 95:30]
  wire [17:0] ___B_2_2_T_5 = $signed(___B_2_2_T_2) + $signed(_B_2_2); // @[calc8x8.scala 95:39]
  wire [17:0] ___B_2_3_T_2 = $signed(_B_2_0) - $signed(_B_2_2); // @[calc8x8.scala 96:30]
  wire [17:0] ___B_2_3_T_5 = $signed(___B_2_3_T_2) - 18'sh0; // @[calc8x8.scala 96:39]
  wire [18:0] ___Bi_2_3_T_3 = {{1{_B_2_1[17]}},_B_2_1}; // @[calc8x8.scala 102:42]
  wire [17:0] ___Bi_2_3_T_5 = ___Bi_2_3_T_3[17:0]; // @[calc8x8.scala 102:42]
  wire [17:0] ___B_3_1_T_2 = $signed(_B_3_0) + $signed(_B_3_1); // @[calc8x8.scala 94:30]
  wire [17:0] ___B_3_1_T_5 = $signed(___B_3_1_T_2) + $signed(_B_3_2); // @[calc8x8.scala 94:39]
  wire [17:0] ___B_3_2_T_2 = $signed(_B_3_0) - $signed(_B_3_1); // @[calc8x8.scala 95:30]
  wire [17:0] ___B_3_2_T_5 = $signed(___B_3_2_T_2) + $signed(_B_3_2); // @[calc8x8.scala 95:39]
  wire [17:0] ___B_3_3_T_2 = $signed(_B_3_0) - $signed(_B_3_2); // @[calc8x8.scala 96:30]
  wire [17:0] ___B_3_3_T_5 = $signed(___B_3_3_T_2) - $signed(_Bi_3_1); // @[calc8x8.scala 96:39]
  wire [17:0] ___B_3_4_T_5 = $signed(___B_3_3_T_2) + $signed(_Bi_3_1); // @[calc8x8.scala 97:39]
  wire [17:0] ___Bi_3_1_T_2 = $signed(_Bi_3_0) + $signed(_Bi_3_1); // @[calc8x8.scala 100:32]
  wire [17:0] ___Bi_3_1_T_5 = $signed(___Bi_3_1_T_2) + $signed(_Bi_3_2); // @[calc8x8.scala 100:42]
  wire [17:0] ___Bi_3_2_T_2 = $signed(_Bi_3_0) - $signed(_Bi_3_1); // @[calc8x8.scala 101:32]
  wire [17:0] ___Bi_3_2_T_5 = $signed(___Bi_3_2_T_2) + $signed(_Bi_3_2); // @[calc8x8.scala 101:42]
  wire [17:0] ___Bi_3_3_T_2 = $signed(_Bi_3_0) - $signed(_Bi_3_2); // @[calc8x8.scala 102:32]
  wire [17:0] ___Bi_3_3_T_5 = $signed(___Bi_3_3_T_2) + $signed(_B_3_1); // @[calc8x8.scala 102:42]
  wire [17:0] ___Bi_3_4_T_5 = $signed(___Bi_3_3_T_2) - $signed(_B_3_1); // @[calc8x8.scala 103:42]
  wire [17:0] ___B_5_1_T_2 = $signed(_B_5_0) + $signed(_B_5_1); // @[calc8x8.scala 94:30]
  wire [17:0] ___B_5_1_T_5 = $signed(___B_5_1_T_2) + $signed(_B_5_2); // @[calc8x8.scala 94:39]
  wire [17:0] ___B_5_2_T_2 = $signed(_B_5_0) - $signed(_B_5_1); // @[calc8x8.scala 95:30]
  wire [17:0] ___B_5_2_T_5 = $signed(___B_5_2_T_2) + $signed(_B_5_2); // @[calc8x8.scala 95:39]
  wire [17:0] ___B_5_3_T_2 = $signed(_B_5_0) - $signed(_B_5_2); // @[calc8x8.scala 96:30]
  wire [17:0] ___B_5_3_T_5 = $signed(___B_5_3_T_2) - 18'sh0; // @[calc8x8.scala 96:39]
  wire [18:0] ___Bi_5_3_T_3 = {{1{_B_5_1[17]}},_B_5_1}; // @[calc8x8.scala 102:42]
  wire [17:0] ___Bi_5_3_T_5 = ___Bi_5_3_T_3[17:0]; // @[calc8x8.scala 102:42]
  wire [18:0] _conv_weight_real_0_T_8 = __B_0_0[18] & ~__B_0_0[17] ? $signed(-19'sh20000) : $signed(__B_0_0); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_0_T_9 = ~__B_0_0[18] & __B_0_0[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_0_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_1_T_8 = __B_0_1[18] & ~__B_0_1[17] ? $signed(-19'sh20000) : $signed(__B_0_1); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_1_T_9 = ~__B_0_1[18] & __B_0_1[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_1_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_2_T_8 = __B_0_2[18] & ~__B_0_2[17] ? $signed(-19'sh20000) : $signed(__B_0_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_2_T_9 = ~__B_0_2[18] & __B_0_2[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_2_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_0_T_2 = $signed(__B_0_3) + $signed(__Bi_0_3); // @[calc8x8.scala 127:59]
  wire [18:0] _conv_weight_comp1_0_T_11 = _conv_weight_comp1_0_T_2[18] & ~_conv_weight_comp1_0_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_0_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_0_T_12 = ~_conv_weight_comp1_0_T_2[18] & _conv_weight_comp1_0_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_0_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_0_T_8 = __B_0_3[18] & ~__B_0_3[17] ? $signed(-19'sh20000) : $signed(__B_0_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_0_T_9 = ~__B_0_3[18] & __B_0_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_0_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_0_T_8 = __Bi_0_3[18] & ~__Bi_0_3[17] ? $signed(-19'sh20000) : $signed(__Bi_0_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_0_T_9 = ~__Bi_0_3[18] & __Bi_0_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_0_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_3_T_8 = __B_0_5[18] & ~__B_0_5[17] ? $signed(-19'sh20000) : $signed(__B_0_5); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_3_T_9 = ~__B_0_5[18] & __B_0_5[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_3_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_4_T_8 = __B_1_0[18] & ~__B_1_0[17] ? $signed(-19'sh20000) : $signed(__B_1_0); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_4_T_9 = ~__B_1_0[18] & __B_1_0[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_4_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_5_T_8 = __B_1_1[18] & ~__B_1_1[17] ? $signed(-19'sh20000) : $signed(__B_1_1); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_5_T_9 = ~__B_1_1[18] & __B_1_1[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_5_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_6_T_8 = __B_1_2[18] & ~__B_1_2[17] ? $signed(-19'sh20000) : $signed(__B_1_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_6_T_9 = ~__B_1_2[18] & __B_1_2[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_6_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_1_T_2 = $signed(__B_1_3) + $signed(__Bi_1_3); // @[calc8x8.scala 127:59]
  wire [18:0] _conv_weight_comp1_1_T_11 = _conv_weight_comp1_1_T_2[18] & ~_conv_weight_comp1_1_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_1_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_1_T_12 = ~_conv_weight_comp1_1_T_2[18] & _conv_weight_comp1_1_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_1_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_1_T_8 = __B_1_3[18] & ~__B_1_3[17] ? $signed(-19'sh20000) : $signed(__B_1_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_1_T_9 = ~__B_1_3[18] & __B_1_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_1_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_1_T_8 = __Bi_1_3[18] & ~__Bi_1_3[17] ? $signed(-19'sh20000) : $signed(__Bi_1_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_1_T_9 = ~__Bi_1_3[18] & __Bi_1_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_1_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_7_T_8 = __B_1_5[18] & ~__B_1_5[17] ? $signed(-19'sh20000) : $signed(__B_1_5); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_7_T_9 = ~__B_1_5[18] & __B_1_5[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_7_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_8_T_8 = __B_2_0[18] & ~__B_2_0[17] ? $signed(-19'sh20000) : $signed(__B_2_0); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_8_T_9 = ~__B_2_0[18] & __B_2_0[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_8_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_9_T_8 = __B_2_1[18] & ~__B_2_1[17] ? $signed(-19'sh20000) : $signed(__B_2_1); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_9_T_9 = ~__B_2_1[18] & __B_2_1[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_9_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_10_T_8 = __B_2_2[18] & ~__B_2_2[17] ? $signed(-19'sh20000) : $signed(__B_2_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_10_T_9 = ~__B_2_2[18] & __B_2_2[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_10_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_2_T_2 = $signed(__B_2_3) + $signed(__Bi_2_3); // @[calc8x8.scala 127:59]
  wire [18:0] _conv_weight_comp1_2_T_11 = _conv_weight_comp1_2_T_2[18] & ~_conv_weight_comp1_2_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_2_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_2_T_12 = ~_conv_weight_comp1_2_T_2[18] & _conv_weight_comp1_2_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_2_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_2_T_8 = __B_2_3[18] & ~__B_2_3[17] ? $signed(-19'sh20000) : $signed(__B_2_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_2_T_9 = ~__B_2_3[18] & __B_2_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_2_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_2_T_8 = __Bi_2_3[18] & ~__Bi_2_3[17] ? $signed(-19'sh20000) : $signed(__Bi_2_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_2_T_9 = ~__Bi_2_3[18] & __Bi_2_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_2_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_11_T_8 = __B_2_5[18] & ~__B_2_5[17] ? $signed(-19'sh20000) : $signed(__B_2_5); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_11_T_9 = ~__B_2_5[18] & __B_2_5[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_11_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_3_T_2 = $signed(__B_3_0) + $signed(__Bi_3_0); // @[calc8x8.scala 122:59]
  wire [18:0] _conv_weight_comp1_3_T_11 = _conv_weight_comp1_3_T_2[18] & ~_conv_weight_comp1_3_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_3_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_3_T_12 = ~_conv_weight_comp1_3_T_2[18] & _conv_weight_comp1_3_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_3_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_3_T_8 = __B_3_0[18] & ~__B_3_0[17] ? $signed(-19'sh20000) : $signed(__B_3_0); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_3_T_9 = ~__B_3_0[18] & __B_3_0[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_3_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_3_T_8 = __Bi_3_0[18] & ~__Bi_3_0[17] ? $signed(-19'sh20000) : $signed(__Bi_3_0); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_3_T_9 = ~__Bi_3_0[18] & __Bi_3_0[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_3_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_4_T_2 = $signed(__B_3_1) + $signed(__Bi_3_1); // @[calc8x8.scala 122:59]
  wire [18:0] _conv_weight_comp1_4_T_11 = _conv_weight_comp1_4_T_2[18] & ~_conv_weight_comp1_4_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_4_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_4_T_12 = ~_conv_weight_comp1_4_T_2[18] & _conv_weight_comp1_4_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_4_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_4_T_8 = __B_3_1[18] & ~__B_3_1[17] ? $signed(-19'sh20000) : $signed(__B_3_1); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_4_T_9 = ~__B_3_1[18] & __B_3_1[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_4_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_4_T_8 = __Bi_3_1[18] & ~__Bi_3_1[17] ? $signed(-19'sh20000) : $signed(__Bi_3_1); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_4_T_9 = ~__Bi_3_1[18] & __Bi_3_1[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_4_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_5_T_2 = $signed(__B_3_2) + $signed(__Bi_3_2); // @[calc8x8.scala 122:59]
  wire [18:0] _conv_weight_comp1_5_T_11 = _conv_weight_comp1_5_T_2[18] & ~_conv_weight_comp1_5_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_5_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_5_T_12 = ~_conv_weight_comp1_5_T_2[18] & _conv_weight_comp1_5_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_5_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_5_T_8 = __B_3_2[18] & ~__B_3_2[17] ? $signed(-19'sh20000) : $signed(__B_3_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_5_T_9 = ~__B_3_2[18] & __B_3_2[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_5_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_5_T_8 = __Bi_3_2[18] & ~__Bi_3_2[17] ? $signed(-19'sh20000) : $signed(__Bi_3_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_5_T_9 = ~__Bi_3_2[18] & __Bi_3_2[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_5_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_6_T_2 = $signed(__B_3_3) + $signed(__Bi_3_3); // @[calc8x8.scala 122:59]
  wire [18:0] _conv_weight_comp1_6_T_11 = _conv_weight_comp1_6_T_2[18] & ~_conv_weight_comp1_6_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_6_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_6_T_12 = ~_conv_weight_comp1_6_T_2[18] & _conv_weight_comp1_6_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_6_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_6_T_8 = __B_3_3[18] & ~__B_3_3[17] ? $signed(-19'sh20000) : $signed(__B_3_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_6_T_9 = ~__B_3_3[18] & __B_3_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_6_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_6_T_8 = __Bi_3_3[18] & ~__Bi_3_3[17] ? $signed(-19'sh20000) : $signed(__Bi_3_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_6_T_9 = ~__Bi_3_3[18] & __Bi_3_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_6_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_7_T_2 = $signed(__B_3_4) + $signed(__Bi_3_4); // @[calc8x8.scala 122:59]
  wire [18:0] _conv_weight_comp1_7_T_11 = _conv_weight_comp1_7_T_2[18] & ~_conv_weight_comp1_7_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_7_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_7_T_12 = ~_conv_weight_comp1_7_T_2[18] & _conv_weight_comp1_7_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_7_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_7_T_8 = __B_3_4[18] & ~__B_3_4[17] ? $signed(-19'sh20000) : $signed(__B_3_4); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_7_T_9 = ~__B_3_4[18] & __B_3_4[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_7_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_7_T_8 = __Bi_3_4[18] & ~__Bi_3_4[17] ? $signed(-19'sh20000) : $signed(__Bi_3_4); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_7_T_9 = ~__Bi_3_4[18] & __Bi_3_4[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_7_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_8_T_2 = $signed(__B_3_5) + $signed(__Bi_3_5); // @[calc8x8.scala 122:59]
  wire [18:0] _conv_weight_comp1_8_T_11 = _conv_weight_comp1_8_T_2[18] & ~_conv_weight_comp1_8_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_8_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_8_T_12 = ~_conv_weight_comp1_8_T_2[18] & _conv_weight_comp1_8_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_8_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_8_T_8 = __B_3_5[18] & ~__B_3_5[17] ? $signed(-19'sh20000) : $signed(__B_3_5); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_8_T_9 = ~__B_3_5[18] & __B_3_5[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_8_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_8_T_8 = __Bi_3_5[18] & ~__Bi_3_5[17] ? $signed(-19'sh20000) : $signed(__Bi_3_5); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_8_T_9 = ~__Bi_3_5[18] & __Bi_3_5[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_8_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_12_T_8 = __B_5_0[18] & ~__B_5_0[17] ? $signed(-19'sh20000) : $signed(__B_5_0); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_12_T_9 = ~__B_5_0[18] & __B_5_0[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_12_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_13_T_8 = __B_5_1[18] & ~__B_5_1[17] ? $signed(-19'sh20000) : $signed(__B_5_1); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_13_T_9 = ~__B_5_1[18] & __B_5_1[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_13_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_14_T_8 = __B_5_2[18] & ~__B_5_2[17] ? $signed(-19'sh20000) : $signed(__B_5_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_14_T_9 = ~__B_5_2[18] & __B_5_2[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_14_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp1_9_T_2 = $signed(__B_5_3) + $signed(__Bi_5_3); // @[calc8x8.scala 127:59]
  wire [18:0] _conv_weight_comp1_9_T_11 = _conv_weight_comp1_9_T_2[18] & ~_conv_weight_comp1_9_T_2[17] ? $signed(-19'sh20000
    ) : $signed(_conv_weight_comp1_9_T_2); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp1_9_T_12 = ~_conv_weight_comp1_9_T_2[18] & _conv_weight_comp1_9_T_2[17] ? $signed(19'sh1ffff
    ) : $signed(_conv_weight_comp1_9_T_11); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp2_9_T_8 = __B_5_3[18] & ~__B_5_3[17] ? $signed(-19'sh20000) : $signed(__B_5_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp2_9_T_9 = ~__B_5_3[18] & __B_5_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp2_9_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_comp3_9_T_8 = __Bi_5_3[18] & ~__Bi_5_3[17] ? $signed(-19'sh20000) : $signed(__Bi_5_3); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_comp3_9_T_9 = ~__Bi_5_3[18] & __Bi_5_3[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_comp3_9_T_8); // @[calc8x8.scala 111:19]
  wire [18:0] _conv_weight_real_15_T_8 = __B_5_5[18] & ~__B_5_5[17] ? $signed(-19'sh20000) : $signed(__B_5_5); // @[calc8x8.scala 111:61]
  wire [18:0] _conv_weight_real_15_T_9 = ~__B_5_5[18] & __B_5_5[17] ? $signed(19'sh1ffff) : $signed(
    _conv_weight_real_15_T_8); // @[calc8x8.scala 111:19]
  wire  _T_2 = 2'h0 == io_flag; // @[Conditional.scala 37:30]
  wire  _T_5 = 2'h1 == io_flag; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h2 == io_flag; // @[Conditional.scala 37:30]
  wire [15:0] _GEN_0 = _T_8 ? $signed(io_input_up_0) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_1 = _T_8 ? $signed(io_input_up_1) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_2 = _T_8 ? $signed(io_input_up_2) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_3 = _T_8 ? $signed(io_input_up_3) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_4 = _T_8 ? $signed(io_input_up_4) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_5 = _T_8 ? $signed(io_input_up_5) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_6 = _T_8 ? $signed(io_input_left_0) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_7 = _T_8 ? $signed(io_input_mat_0) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_8 = _T_8 ? $signed(io_input_mat_1) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_9 = _T_8 ? $signed(io_input_mat_2) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_10 = _T_8 ? $signed(io_input_mat_3) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_11 = _T_8 ? $signed(io_input_mat_4) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_12 = _T_8 ? $signed(io_input_left_1) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_13 = _T_8 ? $signed(io_input_mat_8) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_14 = _T_8 ? $signed(io_input_mat_9) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_15 = _T_8 ? $signed(io_input_mat_10) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_16 = _T_8 ? $signed(io_input_mat_11) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_17 = _T_8 ? $signed(io_input_mat_12) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_18 = _T_8 ? $signed(io_input_left_2) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_19 = _T_8 ? $signed(io_input_mat_16) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_20 = _T_8 ? $signed(io_input_mat_17) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_21 = _T_8 ? $signed(io_input_mat_18) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_22 = _T_8 ? $signed(io_input_mat_19) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_23 = _T_8 ? $signed(io_input_mat_20) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_24 = _T_8 ? $signed(io_input_left_3) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_25 = _T_8 ? $signed(io_input_mat_24) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_26 = _T_8 ? $signed(io_input_mat_25) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_27 = _T_8 ? $signed(io_input_mat_26) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_28 = _T_8 ? $signed(io_input_mat_27) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_29 = _T_8 ? $signed(io_input_mat_28) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_30 = _T_8 ? $signed(io_input_left_4) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_31 = _T_8 ? $signed(io_input_mat_32) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_32 = _T_8 ? $signed(io_input_mat_33) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_33 = _T_8 ? $signed(io_input_mat_34) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_34 = _T_8 ? $signed(io_input_mat_35) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_35 = _T_8 ? $signed(io_input_mat_36) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 163:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_38 = _T_8 ? $signed(io_input_up_6) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_39 = _T_8 ? $signed(io_input_up_7) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_40 = _T_8 ? $signed(io_input_up_8) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_41 = _T_8 ? $signed(io_input_up_9) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_44 = _T_8 ? $signed(io_input_mat_5) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_45 = _T_8 ? $signed(io_input_mat_6) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_46 = _T_8 ? $signed(io_input_mat_7) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_47 = _T_8 ? $signed(io_input_right_0) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_50 = _T_8 ? $signed(io_input_mat_13) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_51 = _T_8 ? $signed(io_input_mat_14) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_52 = _T_8 ? $signed(io_input_mat_15) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_53 = _T_8 ? $signed(io_input_right_1) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_56 = _T_8 ? $signed(io_input_mat_21) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_57 = _T_8 ? $signed(io_input_mat_22) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_58 = _T_8 ? $signed(io_input_mat_23) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_59 = _T_8 ? $signed(io_input_right_2) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_62 = _T_8 ? $signed(io_input_mat_29) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_63 = _T_8 ? $signed(io_input_mat_30) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_64 = _T_8 ? $signed(io_input_mat_31) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_65 = _T_8 ? $signed(io_input_right_3) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_68 = _T_8 ? $signed(io_input_mat_37) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_69 = _T_8 ? $signed(io_input_mat_38) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_70 = _T_8 ? $signed(io_input_mat_39) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_71 = _T_8 ? $signed(io_input_right_4) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 164:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_84 = _T_8 ? $signed(io_input_left_5) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_85 = _T_8 ? $signed(io_input_mat_40) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_86 = _T_8 ? $signed(io_input_mat_41) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_87 = _T_8 ? $signed(io_input_mat_42) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_88 = _T_8 ? $signed(io_input_mat_43) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_89 = _T_8 ? $signed(io_input_mat_44) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_90 = _T_8 ? $signed(io_input_left_6) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_91 = _T_8 ? $signed(io_input_mat_48) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_92 = _T_8 ? $signed(io_input_mat_49) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_93 = _T_8 ? $signed(io_input_mat_50) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_94 = _T_8 ? $signed(io_input_mat_51) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_95 = _T_8 ? $signed(io_input_mat_52) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_96 = _T_8 ? $signed(io_input_left_7) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_97 = _T_8 ? $signed(io_input_mat_56) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_98 = _T_8 ? $signed(io_input_mat_57) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_99 = _T_8 ? $signed(io_input_mat_58) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_100 = _T_8 ? $signed(io_input_mat_59) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_101 = _T_8 ? $signed(io_input_mat_60) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_102 = _T_8 ? $signed(io_input_down_0) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_103 = _T_8 ? $signed(io_input_down_1) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_104 = _T_8 ? $signed(io_input_down_2) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_105 = _T_8 ? $signed(io_input_down_3) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_106 = _T_8 ? $signed(io_input_down_4) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_107 = _T_8 ? $signed(io_input_down_5) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 165:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_122 = _T_8 ? $signed(io_input_mat_45) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_123 = _T_8 ? $signed(io_input_mat_46) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_124 = _T_8 ? $signed(io_input_mat_47) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_125 = _T_8 ? $signed(io_input_right_5) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_128 = _T_8 ? $signed(io_input_mat_53) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_129 = _T_8 ? $signed(io_input_mat_54) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_130 = _T_8 ? $signed(io_input_mat_55) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_131 = _T_8 ? $signed(io_input_right_6) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_134 = _T_8 ? $signed(io_input_mat_61) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_135 = _T_8 ? $signed(io_input_mat_62) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_136 = _T_8 ? $signed(io_input_mat_63) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_137 = _T_8 ? $signed(io_input_right_7) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_140 = _T_8 ? $signed(io_input_down_6) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_141 = _T_8 ? $signed(io_input_down_7) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_142 = _T_8 ? $signed(io_input_down_8) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [15:0] _GEN_143 = _T_8 ? $signed(io_input_down_9) : $signed(16'sh0); // @[Conditional.scala 39:67 calc8x8.scala 166:24 calc8x8.scala 61:20]
  wire [17:0] conv_weight_comp3_0 = _conv_weight_comp3_0_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 129:38]
  wire [17:0] _GEN_144 = _T_8 ? $signed(conv_weight_comp3_0) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_1 = _conv_weight_comp3_1_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 129:38]
  wire [17:0] _GEN_145 = _T_8 ? $signed(conv_weight_comp3_1) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_2 = _conv_weight_comp3_2_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 129:38]
  wire [17:0] _GEN_146 = _T_8 ? $signed(conv_weight_comp3_2) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_3 = _conv_weight_comp3_3_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 124:38]
  wire [17:0] _GEN_147 = _T_8 ? $signed(conv_weight_comp3_3) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_4 = _conv_weight_comp3_4_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 124:38]
  wire [17:0] _GEN_148 = _T_8 ? $signed(conv_weight_comp3_4) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_5 = _conv_weight_comp3_5_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 124:38]
  wire [17:0] _GEN_149 = _T_8 ? $signed(conv_weight_comp3_5) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_6 = _conv_weight_comp3_6_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 124:38]
  wire [17:0] _GEN_150 = _T_8 ? $signed(conv_weight_comp3_6) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_7 = _conv_weight_comp3_7_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 124:38]
  wire [17:0] _GEN_151 = _T_8 ? $signed(conv_weight_comp3_7) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_8 = _conv_weight_comp3_8_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 124:38]
  wire [17:0] _GEN_152 = _T_8 ? $signed(conv_weight_comp3_8) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp3_9 = _conv_weight_comp3_9_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 129:38]
  wire [17:0] _GEN_153 = _T_8 ? $signed(conv_weight_comp3_9) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_0 = _conv_weight_comp2_0_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 128:38]
  wire [17:0] _GEN_154 = _T_8 ? $signed(conv_weight_comp2_0) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_1 = _conv_weight_comp2_1_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 128:38]
  wire [17:0] _GEN_155 = _T_8 ? $signed(conv_weight_comp2_1) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_2 = _conv_weight_comp2_2_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 128:38]
  wire [17:0] _GEN_156 = _T_8 ? $signed(conv_weight_comp2_2) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_3 = _conv_weight_comp2_3_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 123:38]
  wire [17:0] _GEN_157 = _T_8 ? $signed(conv_weight_comp2_3) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_4 = _conv_weight_comp2_4_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 123:38]
  wire [17:0] _GEN_158 = _T_8 ? $signed(conv_weight_comp2_4) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_5 = _conv_weight_comp2_5_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 123:38]
  wire [17:0] _GEN_159 = _T_8 ? $signed(conv_weight_comp2_5) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_6 = _conv_weight_comp2_6_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 123:38]
  wire [17:0] _GEN_160 = _T_8 ? $signed(conv_weight_comp2_6) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_7 = _conv_weight_comp2_7_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 123:38]
  wire [17:0] _GEN_161 = _T_8 ? $signed(conv_weight_comp2_7) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_8 = _conv_weight_comp2_8_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 123:38]
  wire [17:0] _GEN_162 = _T_8 ? $signed(conv_weight_comp2_8) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp2_9 = _conv_weight_comp2_9_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 128:38]
  wire [17:0] _GEN_163 = _T_8 ? $signed(conv_weight_comp2_9) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_0 = _conv_weight_comp1_0_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 127:38]
  wire [17:0] _GEN_164 = _T_8 ? $signed(conv_weight_comp1_0) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_1 = _conv_weight_comp1_1_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 127:38]
  wire [17:0] _GEN_165 = _T_8 ? $signed(conv_weight_comp1_1) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_2 = _conv_weight_comp1_2_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 127:38]
  wire [17:0] _GEN_166 = _T_8 ? $signed(conv_weight_comp1_2) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_3 = _conv_weight_comp1_3_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 122:38]
  wire [17:0] _GEN_167 = _T_8 ? $signed(conv_weight_comp1_3) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_4 = _conv_weight_comp1_4_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 122:38]
  wire [17:0] _GEN_168 = _T_8 ? $signed(conv_weight_comp1_4) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_5 = _conv_weight_comp1_5_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 122:38]
  wire [17:0] _GEN_169 = _T_8 ? $signed(conv_weight_comp1_5) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_6 = _conv_weight_comp1_6_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 122:38]
  wire [17:0] _GEN_170 = _T_8 ? $signed(conv_weight_comp1_6) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_7 = _conv_weight_comp1_7_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 122:38]
  wire [17:0] _GEN_171 = _T_8 ? $signed(conv_weight_comp1_7) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_8 = _conv_weight_comp1_8_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 122:38]
  wire [17:0] _GEN_172 = _T_8 ? $signed(conv_weight_comp1_8) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_comp1_9 = _conv_weight_comp1_9_T_12[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 127:38]
  wire [17:0] _GEN_173 = _T_8 ? $signed(conv_weight_comp1_9) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_0 = _conv_weight_real_0_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_174 = _T_8 ? $signed(conv_weight_real_0) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_1 = _conv_weight_real_1_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_175 = _T_8 ? $signed(conv_weight_real_1) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_2 = _conv_weight_real_2_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_176 = _T_8 ? $signed(conv_weight_real_2) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_3 = _conv_weight_real_3_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_177 = _T_8 ? $signed(conv_weight_real_3) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_4 = _conv_weight_real_4_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_178 = _T_8 ? $signed(conv_weight_real_4) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_5 = _conv_weight_real_5_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_179 = _T_8 ? $signed(conv_weight_real_5) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_6 = _conv_weight_real_6_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_180 = _T_8 ? $signed(conv_weight_real_6) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_7 = _conv_weight_real_7_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_181 = _T_8 ? $signed(conv_weight_real_7) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_8 = _conv_weight_real_8_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_182 = _T_8 ? $signed(conv_weight_real_8) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_9 = _conv_weight_real_9_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_183 = _T_8 ? $signed(conv_weight_real_9) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_10 = _conv_weight_real_10_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_184 = _T_8 ? $signed(conv_weight_real_10) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_11 = _conv_weight_real_11_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_185 = _T_8 ? $signed(conv_weight_real_11) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_12 = _conv_weight_real_12_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_186 = _T_8 ? $signed(conv_weight_real_12) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_13 = _conv_weight_real_13_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_187 = _T_8 ? $signed(conv_weight_real_13) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_14 = _conv_weight_real_14_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_188 = _T_8 ? $signed(conv_weight_real_14) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [17:0] conv_weight_real_15 = _conv_weight_real_15_T_9[17:0]; // @[calc8x8.scala 107:27 calc8x8.scala 119:37]
  wire [17:0] _GEN_189 = _T_8 ? $signed(conv_weight_real_15) : $signed(18'sh0); // @[Conditional.scala 39:67 calc8x8.scala 168:29 calc8x8.scala 63:21]
  wire [1:0] _GEN_190 = _T_8 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 calc8x8.scala 169:27 calc8x8.scala 62:19]
  wire  _GEN_191 = _T_8 & io_valid_in; // @[Conditional.scala 39:67 calc8x8.scala 170:31 calc8x8.scala 64:23]
  wire [36:0] A_0_output_mat_0 = Calc6x6_io_output_mat_0; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_333 = _T_8 ? $signed(A_0_output_mat_0) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_1 = Calc6x6_io_output_mat_1; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_334 = _T_8 ? $signed(A_0_output_mat_1) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_2 = Calc6x6_io_output_mat_2; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_335 = _T_8 ? $signed(A_0_output_mat_2) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_3 = Calc6x6_io_output_mat_3; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_336 = _T_8 ? $signed(A_0_output_mat_3) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_0 = Calc6x6_1_io_output_mat_0; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_337 = _T_8 ? $signed(A_1_output_mat_0) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_1 = Calc6x6_1_io_output_mat_1; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_338 = _T_8 ? $signed(A_1_output_mat_1) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_2 = Calc6x6_1_io_output_mat_2; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_339 = _T_8 ? $signed(A_1_output_mat_2) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_3 = Calc6x6_1_io_output_mat_3; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_340 = _T_8 ? $signed(A_1_output_mat_3) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_4 = Calc6x6_io_output_mat_4; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_341 = _T_8 ? $signed(A_0_output_mat_4) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_5 = Calc6x6_io_output_mat_5; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_342 = _T_8 ? $signed(A_0_output_mat_5) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_6 = Calc6x6_io_output_mat_6; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_343 = _T_8 ? $signed(A_0_output_mat_6) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_7 = Calc6x6_io_output_mat_7; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_344 = _T_8 ? $signed(A_0_output_mat_7) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_4 = Calc6x6_1_io_output_mat_4; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_345 = _T_8 ? $signed(A_1_output_mat_4) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_5 = Calc6x6_1_io_output_mat_5; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_346 = _T_8 ? $signed(A_1_output_mat_5) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_6 = Calc6x6_1_io_output_mat_6; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_347 = _T_8 ? $signed(A_1_output_mat_6) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_7 = Calc6x6_1_io_output_mat_7; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_348 = _T_8 ? $signed(A_1_output_mat_7) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_8 = Calc6x6_io_output_mat_8; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_349 = _T_8 ? $signed(A_0_output_mat_8) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_9 = Calc6x6_io_output_mat_9; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_350 = _T_8 ? $signed(A_0_output_mat_9) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_10 = Calc6x6_io_output_mat_10; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_351 = _T_8 ? $signed(A_0_output_mat_10) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_11 = Calc6x6_io_output_mat_11; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_352 = _T_8 ? $signed(A_0_output_mat_11) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_8 = Calc6x6_1_io_output_mat_8; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_353 = _T_8 ? $signed(A_1_output_mat_8) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_9 = Calc6x6_1_io_output_mat_9; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_354 = _T_8 ? $signed(A_1_output_mat_9) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_10 = Calc6x6_1_io_output_mat_10; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_355 = _T_8 ? $signed(A_1_output_mat_10) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_11 = Calc6x6_1_io_output_mat_11; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_356 = _T_8 ? $signed(A_1_output_mat_11) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_12 = Calc6x6_io_output_mat_12; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_357 = _T_8 ? $signed(A_0_output_mat_12) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_13 = Calc6x6_io_output_mat_13; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_358 = _T_8 ? $signed(A_0_output_mat_13) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_14 = Calc6x6_io_output_mat_14; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_359 = _T_8 ? $signed(A_0_output_mat_14) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_0_output_mat_15 = Calc6x6_io_output_mat_15; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_360 = _T_8 ? $signed(A_0_output_mat_15) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_12 = Calc6x6_1_io_output_mat_12; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_361 = _T_8 ? $signed(A_1_output_mat_12) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_13 = Calc6x6_1_io_output_mat_13; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_362 = _T_8 ? $signed(A_1_output_mat_13) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_14 = Calc6x6_1_io_output_mat_14; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_363 = _T_8 ? $signed(A_1_output_mat_14) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_1_output_mat_15 = Calc6x6_1_io_output_mat_15; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_364 = _T_8 ? $signed(A_1_output_mat_15) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_0 = Calc6x6_2_io_output_mat_0; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_365 = _T_8 ? $signed(A_2_output_mat_0) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_1 = Calc6x6_2_io_output_mat_1; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_366 = _T_8 ? $signed(A_2_output_mat_1) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_2 = Calc6x6_2_io_output_mat_2; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_367 = _T_8 ? $signed(A_2_output_mat_2) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_3 = Calc6x6_2_io_output_mat_3; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_368 = _T_8 ? $signed(A_2_output_mat_3) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_0 = Calc6x6_3_io_output_mat_0; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_369 = _T_8 ? $signed(A_3_output_mat_0) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_1 = Calc6x6_3_io_output_mat_1; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_370 = _T_8 ? $signed(A_3_output_mat_1) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_2 = Calc6x6_3_io_output_mat_2; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_371 = _T_8 ? $signed(A_3_output_mat_2) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_3 = Calc6x6_3_io_output_mat_3; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_372 = _T_8 ? $signed(A_3_output_mat_3) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_4 = Calc6x6_2_io_output_mat_4; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_373 = _T_8 ? $signed(A_2_output_mat_4) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_5 = Calc6x6_2_io_output_mat_5; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_374 = _T_8 ? $signed(A_2_output_mat_5) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_6 = Calc6x6_2_io_output_mat_6; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_375 = _T_8 ? $signed(A_2_output_mat_6) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_7 = Calc6x6_2_io_output_mat_7; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_376 = _T_8 ? $signed(A_2_output_mat_7) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_4 = Calc6x6_3_io_output_mat_4; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_377 = _T_8 ? $signed(A_3_output_mat_4) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_5 = Calc6x6_3_io_output_mat_5; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_378 = _T_8 ? $signed(A_3_output_mat_5) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_6 = Calc6x6_3_io_output_mat_6; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_379 = _T_8 ? $signed(A_3_output_mat_6) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_7 = Calc6x6_3_io_output_mat_7; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_380 = _T_8 ? $signed(A_3_output_mat_7) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_8 = Calc6x6_2_io_output_mat_8; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_381 = _T_8 ? $signed(A_2_output_mat_8) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_9 = Calc6x6_2_io_output_mat_9; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_382 = _T_8 ? $signed(A_2_output_mat_9) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_10 = Calc6x6_2_io_output_mat_10; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_383 = _T_8 ? $signed(A_2_output_mat_10) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_11 = Calc6x6_2_io_output_mat_11; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_384 = _T_8 ? $signed(A_2_output_mat_11) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_8 = Calc6x6_3_io_output_mat_8; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_385 = _T_8 ? $signed(A_3_output_mat_8) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_9 = Calc6x6_3_io_output_mat_9; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_386 = _T_8 ? $signed(A_3_output_mat_9) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_10 = Calc6x6_3_io_output_mat_10; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_387 = _T_8 ? $signed(A_3_output_mat_10) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_11 = Calc6x6_3_io_output_mat_11; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_388 = _T_8 ? $signed(A_3_output_mat_11) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_12 = Calc6x6_2_io_output_mat_12; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_389 = _T_8 ? $signed(A_2_output_mat_12) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_13 = Calc6x6_2_io_output_mat_13; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_390 = _T_8 ? $signed(A_2_output_mat_13) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_14 = Calc6x6_2_io_output_mat_14; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_391 = _T_8 ? $signed(A_2_output_mat_14) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_2_output_mat_15 = Calc6x6_2_io_output_mat_15; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_392 = _T_8 ? $signed(A_2_output_mat_15) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_12 = Calc6x6_3_io_output_mat_12; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_393 = _T_8 ? $signed(A_3_output_mat_12) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_13 = Calc6x6_3_io_output_mat_13; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_394 = _T_8 ? $signed(A_3_output_mat_13) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_14 = Calc6x6_3_io_output_mat_14; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_395 = _T_8 ? $signed(A_3_output_mat_14) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire [36:0] A_3_output_mat_15 = Calc6x6_3_io_output_mat_15; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire [36:0] _GEN_396 = _T_8 ? $signed(A_3_output_mat_15) : $signed(37'sh0); // @[Conditional.scala 39:67 calc8x8.scala 172:23 calc8x8.scala 67:15]
  wire  A_0_valid_out = Calc6x6_io_valid_out; // @[calc8x8.scala 59:20 calc8x8.scala 59:20]
  wire  _GEN_397 = _T_8 & A_0_valid_out; // @[Conditional.scala 39:67 calc8x8.scala 173:26 calc8x8.scala 68:18]
  wire [15:0] _GEN_398 = _T_5 ? $signed(io_input_mat_0) : $signed(_GEN_0); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_399 = _T_5 ? $signed(io_input_mat_1) : $signed(_GEN_1); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_400 = _T_5 ? $signed(io_input_mat_2) : $signed(_GEN_2); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_401 = _T_5 ? $signed(io_input_mat_3) : $signed(_GEN_3); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_402 = _T_5 ? $signed(16'sh0) : $signed(_GEN_4); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_403 = _T_5 ? $signed(16'sh0) : $signed(_GEN_5); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_404 = _T_5 ? $signed(io_input_mat_8) : $signed(_GEN_6); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_405 = _T_5 ? $signed(io_input_mat_9) : $signed(_GEN_7); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_406 = _T_5 ? $signed(io_input_mat_10) : $signed(_GEN_8); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_407 = _T_5 ? $signed(io_input_mat_11) : $signed(_GEN_9); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_408 = _T_5 ? $signed(16'sh0) : $signed(_GEN_10); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_409 = _T_5 ? $signed(16'sh0) : $signed(_GEN_11); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_410 = _T_5 ? $signed(io_input_mat_16) : $signed(_GEN_12); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_411 = _T_5 ? $signed(io_input_mat_17) : $signed(_GEN_13); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_412 = _T_5 ? $signed(io_input_mat_18) : $signed(_GEN_14); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_413 = _T_5 ? $signed(io_input_mat_19) : $signed(_GEN_15); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_414 = _T_5 ? $signed(16'sh0) : $signed(_GEN_16); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_415 = _T_5 ? $signed(16'sh0) : $signed(_GEN_17); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_416 = _T_5 ? $signed(io_input_mat_24) : $signed(_GEN_18); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_417 = _T_5 ? $signed(io_input_mat_25) : $signed(_GEN_19); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_418 = _T_5 ? $signed(io_input_mat_26) : $signed(_GEN_20); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_419 = _T_5 ? $signed(io_input_mat_27) : $signed(_GEN_21); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_420 = _T_5 ? $signed(16'sh0) : $signed(_GEN_22); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_421 = _T_5 ? $signed(16'sh0) : $signed(_GEN_23); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_422 = _T_5 ? $signed(16'sh0) : $signed(_GEN_24); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_423 = _T_5 ? $signed(16'sh0) : $signed(_GEN_25); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_424 = _T_5 ? $signed(16'sh0) : $signed(_GEN_26); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_425 = _T_5 ? $signed(16'sh0) : $signed(_GEN_27); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_426 = _T_5 ? $signed(16'sh0) : $signed(_GEN_28); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_427 = _T_5 ? $signed(16'sh0) : $signed(_GEN_29); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_428 = _T_5 ? $signed(16'sh0) : $signed(_GEN_30); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_429 = _T_5 ? $signed(16'sh0) : $signed(_GEN_31); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_430 = _T_5 ? $signed(16'sh0) : $signed(_GEN_32); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_431 = _T_5 ? $signed(16'sh0) : $signed(_GEN_33); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_432 = _T_5 ? $signed(16'sh0) : $signed(_GEN_34); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_433 = _T_5 ? $signed(16'sh0) : $signed(_GEN_35); // @[Conditional.scala 39:67 calc8x8.scala 150:24]
  wire [15:0] _GEN_434 = _T_5 ? $signed(io_input_mat_3) : $signed(_GEN_4); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_435 = _T_5 ? $signed(io_input_mat_4) : $signed(_GEN_5); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_436 = _T_5 ? $signed(io_input_mat_5) : $signed(_GEN_38); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_437 = _T_5 ? $signed(io_input_mat_6) : $signed(_GEN_39); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_438 = _T_5 ? $signed(io_input_mat_7) : $signed(_GEN_40); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_439 = _T_5 ? $signed(16'sh0) : $signed(_GEN_41); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_440 = _T_5 ? $signed(io_input_mat_11) : $signed(_GEN_10); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_441 = _T_5 ? $signed(io_input_mat_12) : $signed(_GEN_11); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_442 = _T_5 ? $signed(io_input_mat_13) : $signed(_GEN_44); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_443 = _T_5 ? $signed(io_input_mat_14) : $signed(_GEN_45); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_444 = _T_5 ? $signed(io_input_mat_15) : $signed(_GEN_46); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_445 = _T_5 ? $signed(16'sh0) : $signed(_GEN_47); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_446 = _T_5 ? $signed(io_input_mat_19) : $signed(_GEN_16); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_447 = _T_5 ? $signed(io_input_mat_20) : $signed(_GEN_17); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_448 = _T_5 ? $signed(io_input_mat_21) : $signed(_GEN_50); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_449 = _T_5 ? $signed(io_input_mat_22) : $signed(_GEN_51); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_450 = _T_5 ? $signed(io_input_mat_23) : $signed(_GEN_52); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_451 = _T_5 ? $signed(16'sh0) : $signed(_GEN_53); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_452 = _T_5 ? $signed(io_input_mat_27) : $signed(_GEN_22); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_453 = _T_5 ? $signed(io_input_mat_28) : $signed(_GEN_23); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_454 = _T_5 ? $signed(io_input_mat_29) : $signed(_GEN_56); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_455 = _T_5 ? $signed(io_input_mat_30) : $signed(_GEN_57); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_456 = _T_5 ? $signed(io_input_mat_31) : $signed(_GEN_58); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_457 = _T_5 ? $signed(16'sh0) : $signed(_GEN_59); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_460 = _T_5 ? $signed(16'sh0) : $signed(_GEN_62); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_461 = _T_5 ? $signed(16'sh0) : $signed(_GEN_63); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_462 = _T_5 ? $signed(16'sh0) : $signed(_GEN_64); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_463 = _T_5 ? $signed(16'sh0) : $signed(_GEN_65); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_466 = _T_5 ? $signed(16'sh0) : $signed(_GEN_68); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_467 = _T_5 ? $signed(16'sh0) : $signed(_GEN_69); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_468 = _T_5 ? $signed(16'sh0) : $signed(_GEN_70); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_469 = _T_5 ? $signed(16'sh0) : $signed(_GEN_71); // @[Conditional.scala 39:67 calc8x8.scala 151:24]
  wire [15:0] _GEN_470 = _T_5 ? $signed(io_input_mat_24) : $signed(_GEN_24); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_471 = _T_5 ? $signed(io_input_mat_25) : $signed(_GEN_25); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_472 = _T_5 ? $signed(io_input_mat_26) : $signed(_GEN_26); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_473 = _T_5 ? $signed(io_input_mat_27) : $signed(_GEN_27); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_476 = _T_5 ? $signed(io_input_mat_32) : $signed(_GEN_30); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_477 = _T_5 ? $signed(io_input_mat_33) : $signed(_GEN_31); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_478 = _T_5 ? $signed(io_input_mat_34) : $signed(_GEN_32); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_479 = _T_5 ? $signed(io_input_mat_35) : $signed(_GEN_33); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_482 = _T_5 ? $signed(io_input_mat_40) : $signed(_GEN_84); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_483 = _T_5 ? $signed(io_input_mat_41) : $signed(_GEN_85); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_484 = _T_5 ? $signed(io_input_mat_42) : $signed(_GEN_86); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_485 = _T_5 ? $signed(io_input_mat_43) : $signed(_GEN_87); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_486 = _T_5 ? $signed(16'sh0) : $signed(_GEN_88); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_487 = _T_5 ? $signed(16'sh0) : $signed(_GEN_89); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_488 = _T_5 ? $signed(io_input_mat_48) : $signed(_GEN_90); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_489 = _T_5 ? $signed(io_input_mat_49) : $signed(_GEN_91); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_490 = _T_5 ? $signed(io_input_mat_50) : $signed(_GEN_92); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_491 = _T_5 ? $signed(io_input_mat_51) : $signed(_GEN_93); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_492 = _T_5 ? $signed(16'sh0) : $signed(_GEN_94); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_493 = _T_5 ? $signed(16'sh0) : $signed(_GEN_95); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_494 = _T_5 ? $signed(io_input_mat_56) : $signed(_GEN_96); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_495 = _T_5 ? $signed(io_input_mat_57) : $signed(_GEN_97); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_496 = _T_5 ? $signed(io_input_mat_58) : $signed(_GEN_98); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_497 = _T_5 ? $signed(io_input_mat_59) : $signed(_GEN_99); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_498 = _T_5 ? $signed(16'sh0) : $signed(_GEN_100); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_499 = _T_5 ? $signed(16'sh0) : $signed(_GEN_101); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_500 = _T_5 ? $signed(16'sh0) : $signed(_GEN_102); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_501 = _T_5 ? $signed(16'sh0) : $signed(_GEN_103); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_502 = _T_5 ? $signed(16'sh0) : $signed(_GEN_104); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_503 = _T_5 ? $signed(16'sh0) : $signed(_GEN_105); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_504 = _T_5 ? $signed(16'sh0) : $signed(_GEN_106); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_505 = _T_5 ? $signed(16'sh0) : $signed(_GEN_107); // @[Conditional.scala 39:67 calc8x8.scala 152:24]
  wire [15:0] _GEN_506 = _T_5 ? $signed(io_input_mat_27) : $signed(_GEN_28); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_507 = _T_5 ? $signed(io_input_mat_28) : $signed(_GEN_29); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_508 = _T_5 ? $signed(io_input_mat_29) : $signed(_GEN_62); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_509 = _T_5 ? $signed(io_input_mat_30) : $signed(_GEN_63); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_510 = _T_5 ? $signed(io_input_mat_31) : $signed(_GEN_64); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_512 = _T_5 ? $signed(io_input_mat_35) : $signed(_GEN_34); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_513 = _T_5 ? $signed(io_input_mat_36) : $signed(_GEN_35); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_514 = _T_5 ? $signed(io_input_mat_37) : $signed(_GEN_68); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_515 = _T_5 ? $signed(io_input_mat_38) : $signed(_GEN_69); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_516 = _T_5 ? $signed(io_input_mat_39) : $signed(_GEN_70); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_518 = _T_5 ? $signed(io_input_mat_43) : $signed(_GEN_88); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_519 = _T_5 ? $signed(io_input_mat_44) : $signed(_GEN_89); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_520 = _T_5 ? $signed(io_input_mat_45) : $signed(_GEN_122); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_521 = _T_5 ? $signed(io_input_mat_46) : $signed(_GEN_123); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_522 = _T_5 ? $signed(io_input_mat_47) : $signed(_GEN_124); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_523 = _T_5 ? $signed(16'sh0) : $signed(_GEN_125); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_524 = _T_5 ? $signed(io_input_mat_51) : $signed(_GEN_94); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_525 = _T_5 ? $signed(io_input_mat_52) : $signed(_GEN_95); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_526 = _T_5 ? $signed(io_input_mat_53) : $signed(_GEN_128); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_527 = _T_5 ? $signed(io_input_mat_54) : $signed(_GEN_129); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_528 = _T_5 ? $signed(io_input_mat_55) : $signed(_GEN_130); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_529 = _T_5 ? $signed(16'sh0) : $signed(_GEN_131); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_530 = _T_5 ? $signed(io_input_mat_59) : $signed(_GEN_100); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_531 = _T_5 ? $signed(io_input_mat_60) : $signed(_GEN_101); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_532 = _T_5 ? $signed(io_input_mat_61) : $signed(_GEN_134); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_533 = _T_5 ? $signed(io_input_mat_62) : $signed(_GEN_135); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_534 = _T_5 ? $signed(io_input_mat_63) : $signed(_GEN_136); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_535 = _T_5 ? $signed(16'sh0) : $signed(_GEN_137); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_538 = _T_5 ? $signed(16'sh0) : $signed(_GEN_140); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_539 = _T_5 ? $signed(16'sh0) : $signed(_GEN_141); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_540 = _T_5 ? $signed(16'sh0) : $signed(_GEN_142); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [15:0] _GEN_541 = _T_5 ? $signed(16'sh0) : $signed(_GEN_143); // @[Conditional.scala 39:67 calc8x8.scala 153:24]
  wire [17:0] _GEN_542 = _T_5 ? $signed({{2{io_weight_0_real_0[15]}},io_weight_0_real_0}) : $signed(_GEN_174); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_543 = _T_5 ? $signed({{2{io_weight_0_real_1[15]}},io_weight_0_real_1}) : $signed(_GEN_175); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_544 = _T_5 ? $signed({{2{io_weight_0_real_2[15]}},io_weight_0_real_2}) : $signed(_GEN_176); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_545 = _T_5 ? $signed({{2{io_weight_0_real_3[15]}},io_weight_0_real_3}) : $signed(_GEN_177); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_546 = _T_5 ? $signed({{2{io_weight_0_real_4[15]}},io_weight_0_real_4}) : $signed(_GEN_178); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_547 = _T_5 ? $signed({{2{io_weight_0_real_5[15]}},io_weight_0_real_5}) : $signed(_GEN_179); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_548 = _T_5 ? $signed({{2{io_weight_0_real_6[15]}},io_weight_0_real_6}) : $signed(_GEN_180); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_549 = _T_5 ? $signed({{2{io_weight_0_real_7[15]}},io_weight_0_real_7}) : $signed(_GEN_181); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_550 = _T_5 ? $signed({{2{io_weight_0_real_8[15]}},io_weight_0_real_8}) : $signed(_GEN_182); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_551 = _T_5 ? $signed({{2{io_weight_0_real_9[15]}},io_weight_0_real_9}) : $signed(_GEN_183); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_552 = _T_5 ? $signed({{2{io_weight_0_real_10[15]}},io_weight_0_real_10}) : $signed(_GEN_184); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_553 = _T_5 ? $signed({{2{io_weight_0_real_11[15]}},io_weight_0_real_11}) : $signed(_GEN_185); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_554 = _T_5 ? $signed({{2{io_weight_0_real_12[15]}},io_weight_0_real_12}) : $signed(_GEN_186); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_555 = _T_5 ? $signed({{2{io_weight_0_real_13[15]}},io_weight_0_real_13}) : $signed(_GEN_187); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_556 = _T_5 ? $signed({{2{io_weight_0_real_14[15]}},io_weight_0_real_14}) : $signed(_GEN_188); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_557 = _T_5 ? $signed({{2{io_weight_0_real_15[15]}},io_weight_0_real_15}) : $signed(_GEN_189); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [1:0] _GEN_558 = _T_5 ? 2'h1 : _GEN_190; // @[Conditional.scala 39:67 calc8x8.scala 156:27]
  wire  _GEN_559 = _T_5 ? io_valid_in : _GEN_191; // @[Conditional.scala 39:67 calc8x8.scala 157:31]
  wire [17:0] _GEN_560 = _T_5 ? $signed({{2{io_weight_1_real_0[15]}},io_weight_1_real_0}) : $signed(_GEN_174); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_561 = _T_5 ? $signed({{2{io_weight_1_real_1[15]}},io_weight_1_real_1}) : $signed(_GEN_175); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_562 = _T_5 ? $signed({{2{io_weight_1_real_2[15]}},io_weight_1_real_2}) : $signed(_GEN_176); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_563 = _T_5 ? $signed({{2{io_weight_1_real_3[15]}},io_weight_1_real_3}) : $signed(_GEN_177); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_564 = _T_5 ? $signed({{2{io_weight_1_real_4[15]}},io_weight_1_real_4}) : $signed(_GEN_178); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_565 = _T_5 ? $signed({{2{io_weight_1_real_5[15]}},io_weight_1_real_5}) : $signed(_GEN_179); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_566 = _T_5 ? $signed({{2{io_weight_1_real_6[15]}},io_weight_1_real_6}) : $signed(_GEN_180); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_567 = _T_5 ? $signed({{2{io_weight_1_real_7[15]}},io_weight_1_real_7}) : $signed(_GEN_181); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_568 = _T_5 ? $signed({{2{io_weight_1_real_8[15]}},io_weight_1_real_8}) : $signed(_GEN_182); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_569 = _T_5 ? $signed({{2{io_weight_1_real_9[15]}},io_weight_1_real_9}) : $signed(_GEN_183); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_570 = _T_5 ? $signed({{2{io_weight_1_real_10[15]}},io_weight_1_real_10}) : $signed(_GEN_184); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_571 = _T_5 ? $signed({{2{io_weight_1_real_11[15]}},io_weight_1_real_11}) : $signed(_GEN_185); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_572 = _T_5 ? $signed({{2{io_weight_1_real_12[15]}},io_weight_1_real_12}) : $signed(_GEN_186); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_573 = _T_5 ? $signed({{2{io_weight_1_real_13[15]}},io_weight_1_real_13}) : $signed(_GEN_187); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_574 = _T_5 ? $signed({{2{io_weight_1_real_14[15]}},io_weight_1_real_14}) : $signed(_GEN_188); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_575 = _T_5 ? $signed({{2{io_weight_1_real_15[15]}},io_weight_1_real_15}) : $signed(_GEN_189); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_577 = _T_5 ? $signed({{2{io_weight_2_real_0[15]}},io_weight_2_real_0}) : $signed(_GEN_174); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_578 = _T_5 ? $signed({{2{io_weight_2_real_1[15]}},io_weight_2_real_1}) : $signed(_GEN_175); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_579 = _T_5 ? $signed({{2{io_weight_2_real_2[15]}},io_weight_2_real_2}) : $signed(_GEN_176); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_580 = _T_5 ? $signed({{2{io_weight_2_real_3[15]}},io_weight_2_real_3}) : $signed(_GEN_177); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_581 = _T_5 ? $signed({{2{io_weight_2_real_4[15]}},io_weight_2_real_4}) : $signed(_GEN_178); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_582 = _T_5 ? $signed({{2{io_weight_2_real_5[15]}},io_weight_2_real_5}) : $signed(_GEN_179); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_583 = _T_5 ? $signed({{2{io_weight_2_real_6[15]}},io_weight_2_real_6}) : $signed(_GEN_180); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_584 = _T_5 ? $signed({{2{io_weight_2_real_7[15]}},io_weight_2_real_7}) : $signed(_GEN_181); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_585 = _T_5 ? $signed({{2{io_weight_2_real_8[15]}},io_weight_2_real_8}) : $signed(_GEN_182); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_586 = _T_5 ? $signed({{2{io_weight_2_real_9[15]}},io_weight_2_real_9}) : $signed(_GEN_183); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_587 = _T_5 ? $signed({{2{io_weight_2_real_10[15]}},io_weight_2_real_10}) : $signed(_GEN_184); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_588 = _T_5 ? $signed({{2{io_weight_2_real_11[15]}},io_weight_2_real_11}) : $signed(_GEN_185); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_589 = _T_5 ? $signed({{2{io_weight_2_real_12[15]}},io_weight_2_real_12}) : $signed(_GEN_186); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_590 = _T_5 ? $signed({{2{io_weight_2_real_13[15]}},io_weight_2_real_13}) : $signed(_GEN_187); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_591 = _T_5 ? $signed({{2{io_weight_2_real_14[15]}},io_weight_2_real_14}) : $signed(_GEN_188); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_592 = _T_5 ? $signed({{2{io_weight_2_real_15[15]}},io_weight_2_real_15}) : $signed(_GEN_189); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_594 = _T_5 ? $signed({{2{io_weight_3_real_0[15]}},io_weight_3_real_0}) : $signed(_GEN_174); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_595 = _T_5 ? $signed({{2{io_weight_3_real_1[15]}},io_weight_3_real_1}) : $signed(_GEN_175); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_596 = _T_5 ? $signed({{2{io_weight_3_real_2[15]}},io_weight_3_real_2}) : $signed(_GEN_176); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_597 = _T_5 ? $signed({{2{io_weight_3_real_3[15]}},io_weight_3_real_3}) : $signed(_GEN_177); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_598 = _T_5 ? $signed({{2{io_weight_3_real_4[15]}},io_weight_3_real_4}) : $signed(_GEN_178); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_599 = _T_5 ? $signed({{2{io_weight_3_real_5[15]}},io_weight_3_real_5}) : $signed(_GEN_179); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_600 = _T_5 ? $signed({{2{io_weight_3_real_6[15]}},io_weight_3_real_6}) : $signed(_GEN_180); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_601 = _T_5 ? $signed({{2{io_weight_3_real_7[15]}},io_weight_3_real_7}) : $signed(_GEN_181); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_602 = _T_5 ? $signed({{2{io_weight_3_real_8[15]}},io_weight_3_real_8}) : $signed(_GEN_182); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_603 = _T_5 ? $signed({{2{io_weight_3_real_9[15]}},io_weight_3_real_9}) : $signed(_GEN_183); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_604 = _T_5 ? $signed({{2{io_weight_3_real_10[15]}},io_weight_3_real_10}) : $signed(_GEN_184); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_605 = _T_5 ? $signed({{2{io_weight_3_real_11[15]}},io_weight_3_real_11}) : $signed(_GEN_185); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_606 = _T_5 ? $signed({{2{io_weight_3_real_12[15]}},io_weight_3_real_12}) : $signed(_GEN_186); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_607 = _T_5 ? $signed({{2{io_weight_3_real_13[15]}},io_weight_3_real_13}) : $signed(_GEN_187); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_608 = _T_5 ? $signed({{2{io_weight_3_real_14[15]}},io_weight_3_real_14}) : $signed(_GEN_188); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [17:0] _GEN_609 = _T_5 ? $signed({{2{io_weight_3_real_15[15]}},io_weight_3_real_15}) : $signed(_GEN_189); // @[Conditional.scala 39:67 calc8x8.scala 155:34]
  wire [36:0] _GEN_611 = _T_5 ? $signed(A_0_output_mat_0) : $signed(_GEN_333); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_612 = _T_5 ? $signed(A_0_output_mat_1) : $signed(_GEN_334); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_613 = _T_5 ? $signed(A_0_output_mat_2) : $signed(_GEN_335); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_614 = _T_5 ? $signed(A_0_output_mat_3) : $signed(_GEN_336); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_615 = _T_5 ? $signed(A_1_output_mat_0) : $signed(_GEN_337); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_616 = _T_5 ? $signed(A_1_output_mat_1) : $signed(_GEN_338); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_617 = _T_5 ? $signed(A_1_output_mat_2) : $signed(_GEN_339); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_618 = _T_5 ? $signed(A_1_output_mat_3) : $signed(_GEN_340); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_619 = _T_5 ? $signed(A_0_output_mat_4) : $signed(_GEN_341); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_620 = _T_5 ? $signed(A_0_output_mat_5) : $signed(_GEN_342); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_621 = _T_5 ? $signed(A_0_output_mat_6) : $signed(_GEN_343); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_622 = _T_5 ? $signed(A_0_output_mat_7) : $signed(_GEN_344); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_623 = _T_5 ? $signed(A_1_output_mat_4) : $signed(_GEN_345); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_624 = _T_5 ? $signed(A_1_output_mat_5) : $signed(_GEN_346); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_625 = _T_5 ? $signed(A_1_output_mat_6) : $signed(_GEN_347); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_626 = _T_5 ? $signed(A_1_output_mat_7) : $signed(_GEN_348); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_627 = _T_5 ? $signed(A_0_output_mat_8) : $signed(_GEN_349); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_628 = _T_5 ? $signed(A_0_output_mat_9) : $signed(_GEN_350); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_629 = _T_5 ? $signed(A_0_output_mat_10) : $signed(_GEN_351); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_630 = _T_5 ? $signed(A_0_output_mat_11) : $signed(_GEN_352); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_631 = _T_5 ? $signed(A_1_output_mat_8) : $signed(_GEN_353); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_632 = _T_5 ? $signed(A_1_output_mat_9) : $signed(_GEN_354); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_633 = _T_5 ? $signed(A_1_output_mat_10) : $signed(_GEN_355); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_634 = _T_5 ? $signed(A_1_output_mat_11) : $signed(_GEN_356); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_635 = _T_5 ? $signed(A_0_output_mat_12) : $signed(_GEN_357); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_636 = _T_5 ? $signed(A_0_output_mat_13) : $signed(_GEN_358); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_637 = _T_5 ? $signed(A_0_output_mat_14) : $signed(_GEN_359); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_638 = _T_5 ? $signed(A_0_output_mat_15) : $signed(_GEN_360); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_639 = _T_5 ? $signed(A_1_output_mat_12) : $signed(_GEN_361); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_640 = _T_5 ? $signed(A_1_output_mat_13) : $signed(_GEN_362); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_641 = _T_5 ? $signed(A_1_output_mat_14) : $signed(_GEN_363); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_642 = _T_5 ? $signed(A_1_output_mat_15) : $signed(_GEN_364); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_643 = _T_5 ? $signed(A_2_output_mat_0) : $signed(_GEN_365); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_644 = _T_5 ? $signed(A_2_output_mat_1) : $signed(_GEN_366); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_645 = _T_5 ? $signed(A_2_output_mat_2) : $signed(_GEN_367); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_646 = _T_5 ? $signed(A_2_output_mat_3) : $signed(_GEN_368); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_647 = _T_5 ? $signed(A_3_output_mat_0) : $signed(_GEN_369); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_648 = _T_5 ? $signed(A_3_output_mat_1) : $signed(_GEN_370); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_649 = _T_5 ? $signed(A_3_output_mat_2) : $signed(_GEN_371); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_650 = _T_5 ? $signed(A_3_output_mat_3) : $signed(_GEN_372); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_651 = _T_5 ? $signed(A_2_output_mat_4) : $signed(_GEN_373); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_652 = _T_5 ? $signed(A_2_output_mat_5) : $signed(_GEN_374); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_653 = _T_5 ? $signed(A_2_output_mat_6) : $signed(_GEN_375); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_654 = _T_5 ? $signed(A_2_output_mat_7) : $signed(_GEN_376); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_655 = _T_5 ? $signed(A_3_output_mat_4) : $signed(_GEN_377); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_656 = _T_5 ? $signed(A_3_output_mat_5) : $signed(_GEN_378); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_657 = _T_5 ? $signed(A_3_output_mat_6) : $signed(_GEN_379); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_658 = _T_5 ? $signed(A_3_output_mat_7) : $signed(_GEN_380); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_659 = _T_5 ? $signed(A_2_output_mat_8) : $signed(_GEN_381); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_660 = _T_5 ? $signed(A_2_output_mat_9) : $signed(_GEN_382); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_661 = _T_5 ? $signed(A_2_output_mat_10) : $signed(_GEN_383); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_662 = _T_5 ? $signed(A_2_output_mat_11) : $signed(_GEN_384); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_663 = _T_5 ? $signed(A_3_output_mat_8) : $signed(_GEN_385); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_664 = _T_5 ? $signed(A_3_output_mat_9) : $signed(_GEN_386); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_665 = _T_5 ? $signed(A_3_output_mat_10) : $signed(_GEN_387); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_666 = _T_5 ? $signed(A_3_output_mat_11) : $signed(_GEN_388); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_667 = _T_5 ? $signed(A_2_output_mat_12) : $signed(_GEN_389); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_668 = _T_5 ? $signed(A_2_output_mat_13) : $signed(_GEN_390); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_669 = _T_5 ? $signed(A_2_output_mat_14) : $signed(_GEN_391); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_670 = _T_5 ? $signed(A_2_output_mat_15) : $signed(_GEN_392); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_671 = _T_5 ? $signed(A_3_output_mat_12) : $signed(_GEN_393); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_672 = _T_5 ? $signed(A_3_output_mat_13) : $signed(_GEN_394); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_673 = _T_5 ? $signed(A_3_output_mat_14) : $signed(_GEN_395); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire [36:0] _GEN_674 = _T_5 ? $signed(A_3_output_mat_15) : $signed(_GEN_396); // @[Conditional.scala 39:67 calc8x8.scala 159:23]
  wire  _GEN_675 = _T_5 ? A_0_valid_out : _GEN_397; // @[Conditional.scala 39:67 calc8x8.scala 160:26]
  wire [17:0] _GEN_676 = _T_5 ? $signed(18'sh0) : $signed(_GEN_144); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_677 = _T_5 ? $signed(18'sh0) : $signed(_GEN_145); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_678 = _T_5 ? $signed(18'sh0) : $signed(_GEN_146); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_679 = _T_5 ? $signed(18'sh0) : $signed(_GEN_147); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_680 = _T_5 ? $signed(18'sh0) : $signed(_GEN_148); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_681 = _T_5 ? $signed(18'sh0) : $signed(_GEN_149); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_682 = _T_5 ? $signed(18'sh0) : $signed(_GEN_150); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_683 = _T_5 ? $signed(18'sh0) : $signed(_GEN_151); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_684 = _T_5 ? $signed(18'sh0) : $signed(_GEN_152); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_685 = _T_5 ? $signed(18'sh0) : $signed(_GEN_153); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_686 = _T_5 ? $signed(18'sh0) : $signed(_GEN_154); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_687 = _T_5 ? $signed(18'sh0) : $signed(_GEN_155); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_688 = _T_5 ? $signed(18'sh0) : $signed(_GEN_156); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_689 = _T_5 ? $signed(18'sh0) : $signed(_GEN_157); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_690 = _T_5 ? $signed(18'sh0) : $signed(_GEN_158); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_691 = _T_5 ? $signed(18'sh0) : $signed(_GEN_159); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_692 = _T_5 ? $signed(18'sh0) : $signed(_GEN_160); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_693 = _T_5 ? $signed(18'sh0) : $signed(_GEN_161); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_694 = _T_5 ? $signed(18'sh0) : $signed(_GEN_162); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_695 = _T_5 ? $signed(18'sh0) : $signed(_GEN_163); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_696 = _T_5 ? $signed(18'sh0) : $signed(_GEN_164); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_697 = _T_5 ? $signed(18'sh0) : $signed(_GEN_165); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_698 = _T_5 ? $signed(18'sh0) : $signed(_GEN_166); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_699 = _T_5 ? $signed(18'sh0) : $signed(_GEN_167); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_700 = _T_5 ? $signed(18'sh0) : $signed(_GEN_168); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_701 = _T_5 ? $signed(18'sh0) : $signed(_GEN_169); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_702 = _T_5 ? $signed(18'sh0) : $signed(_GEN_170); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_703 = _T_5 ? $signed(18'sh0) : $signed(_GEN_171); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_704 = _T_5 ? $signed(18'sh0) : $signed(_GEN_172); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  wire [17:0] _GEN_705 = _T_5 ? $signed(18'sh0) : $signed(_GEN_173); // @[Conditional.scala 39:67 calc8x8.scala 63:21]
  Calc6x6 Calc6x6 ( // @[calc8x8.scala 59:39]
    .clock(Calc6x6_clock),
    .reset(Calc6x6_reset),
    .io_input_mat_0(Calc6x6_io_input_mat_0),
    .io_input_mat_1(Calc6x6_io_input_mat_1),
    .io_input_mat_2(Calc6x6_io_input_mat_2),
    .io_input_mat_3(Calc6x6_io_input_mat_3),
    .io_input_mat_4(Calc6x6_io_input_mat_4),
    .io_input_mat_5(Calc6x6_io_input_mat_5),
    .io_input_mat_6(Calc6x6_io_input_mat_6),
    .io_input_mat_7(Calc6x6_io_input_mat_7),
    .io_input_mat_8(Calc6x6_io_input_mat_8),
    .io_input_mat_9(Calc6x6_io_input_mat_9),
    .io_input_mat_10(Calc6x6_io_input_mat_10),
    .io_input_mat_11(Calc6x6_io_input_mat_11),
    .io_input_mat_12(Calc6x6_io_input_mat_12),
    .io_input_mat_13(Calc6x6_io_input_mat_13),
    .io_input_mat_14(Calc6x6_io_input_mat_14),
    .io_input_mat_15(Calc6x6_io_input_mat_15),
    .io_input_mat_16(Calc6x6_io_input_mat_16),
    .io_input_mat_17(Calc6x6_io_input_mat_17),
    .io_input_mat_18(Calc6x6_io_input_mat_18),
    .io_input_mat_19(Calc6x6_io_input_mat_19),
    .io_input_mat_20(Calc6x6_io_input_mat_20),
    .io_input_mat_21(Calc6x6_io_input_mat_21),
    .io_input_mat_22(Calc6x6_io_input_mat_22),
    .io_input_mat_23(Calc6x6_io_input_mat_23),
    .io_input_mat_24(Calc6x6_io_input_mat_24),
    .io_input_mat_25(Calc6x6_io_input_mat_25),
    .io_input_mat_26(Calc6x6_io_input_mat_26),
    .io_input_mat_27(Calc6x6_io_input_mat_27),
    .io_input_mat_28(Calc6x6_io_input_mat_28),
    .io_input_mat_29(Calc6x6_io_input_mat_29),
    .io_input_mat_30(Calc6x6_io_input_mat_30),
    .io_input_mat_31(Calc6x6_io_input_mat_31),
    .io_input_mat_32(Calc6x6_io_input_mat_32),
    .io_input_mat_33(Calc6x6_io_input_mat_33),
    .io_input_mat_34(Calc6x6_io_input_mat_34),
    .io_input_mat_35(Calc6x6_io_input_mat_35),
    .io_flag(Calc6x6_io_flag),
    .io_weight_real_0(Calc6x6_io_weight_real_0),
    .io_weight_real_1(Calc6x6_io_weight_real_1),
    .io_weight_real_2(Calc6x6_io_weight_real_2),
    .io_weight_real_3(Calc6x6_io_weight_real_3),
    .io_weight_real_4(Calc6x6_io_weight_real_4),
    .io_weight_real_5(Calc6x6_io_weight_real_5),
    .io_weight_real_6(Calc6x6_io_weight_real_6),
    .io_weight_real_7(Calc6x6_io_weight_real_7),
    .io_weight_real_8(Calc6x6_io_weight_real_8),
    .io_weight_real_9(Calc6x6_io_weight_real_9),
    .io_weight_real_10(Calc6x6_io_weight_real_10),
    .io_weight_real_11(Calc6x6_io_weight_real_11),
    .io_weight_real_12(Calc6x6_io_weight_real_12),
    .io_weight_real_13(Calc6x6_io_weight_real_13),
    .io_weight_real_14(Calc6x6_io_weight_real_14),
    .io_weight_real_15(Calc6x6_io_weight_real_15),
    .io_weight_comp1_0(Calc6x6_io_weight_comp1_0),
    .io_weight_comp1_1(Calc6x6_io_weight_comp1_1),
    .io_weight_comp1_2(Calc6x6_io_weight_comp1_2),
    .io_weight_comp1_3(Calc6x6_io_weight_comp1_3),
    .io_weight_comp1_4(Calc6x6_io_weight_comp1_4),
    .io_weight_comp1_5(Calc6x6_io_weight_comp1_5),
    .io_weight_comp1_6(Calc6x6_io_weight_comp1_6),
    .io_weight_comp1_7(Calc6x6_io_weight_comp1_7),
    .io_weight_comp1_8(Calc6x6_io_weight_comp1_8),
    .io_weight_comp1_9(Calc6x6_io_weight_comp1_9),
    .io_weight_comp2_0(Calc6x6_io_weight_comp2_0),
    .io_weight_comp2_1(Calc6x6_io_weight_comp2_1),
    .io_weight_comp2_2(Calc6x6_io_weight_comp2_2),
    .io_weight_comp2_3(Calc6x6_io_weight_comp2_3),
    .io_weight_comp2_4(Calc6x6_io_weight_comp2_4),
    .io_weight_comp2_5(Calc6x6_io_weight_comp2_5),
    .io_weight_comp2_6(Calc6x6_io_weight_comp2_6),
    .io_weight_comp2_7(Calc6x6_io_weight_comp2_7),
    .io_weight_comp2_8(Calc6x6_io_weight_comp2_8),
    .io_weight_comp2_9(Calc6x6_io_weight_comp2_9),
    .io_weight_comp3_0(Calc6x6_io_weight_comp3_0),
    .io_weight_comp3_1(Calc6x6_io_weight_comp3_1),
    .io_weight_comp3_2(Calc6x6_io_weight_comp3_2),
    .io_weight_comp3_3(Calc6x6_io_weight_comp3_3),
    .io_weight_comp3_4(Calc6x6_io_weight_comp3_4),
    .io_weight_comp3_5(Calc6x6_io_weight_comp3_5),
    .io_weight_comp3_6(Calc6x6_io_weight_comp3_6),
    .io_weight_comp3_7(Calc6x6_io_weight_comp3_7),
    .io_weight_comp3_8(Calc6x6_io_weight_comp3_8),
    .io_weight_comp3_9(Calc6x6_io_weight_comp3_9),
    .io_output_mat_0(Calc6x6_io_output_mat_0),
    .io_output_mat_1(Calc6x6_io_output_mat_1),
    .io_output_mat_2(Calc6x6_io_output_mat_2),
    .io_output_mat_3(Calc6x6_io_output_mat_3),
    .io_output_mat_4(Calc6x6_io_output_mat_4),
    .io_output_mat_5(Calc6x6_io_output_mat_5),
    .io_output_mat_6(Calc6x6_io_output_mat_6),
    .io_output_mat_7(Calc6x6_io_output_mat_7),
    .io_output_mat_8(Calc6x6_io_output_mat_8),
    .io_output_mat_9(Calc6x6_io_output_mat_9),
    .io_output_mat_10(Calc6x6_io_output_mat_10),
    .io_output_mat_11(Calc6x6_io_output_mat_11),
    .io_output_mat_12(Calc6x6_io_output_mat_12),
    .io_output_mat_13(Calc6x6_io_output_mat_13),
    .io_output_mat_14(Calc6x6_io_output_mat_14),
    .io_output_mat_15(Calc6x6_io_output_mat_15),
    .io_valid_in(Calc6x6_io_valid_in),
    .io_valid_out(Calc6x6_io_valid_out)
  );
  Calc6x6 Calc6x6_1 ( // @[calc8x8.scala 59:39]
    .clock(Calc6x6_1_clock),
    .reset(Calc6x6_1_reset),
    .io_input_mat_0(Calc6x6_1_io_input_mat_0),
    .io_input_mat_1(Calc6x6_1_io_input_mat_1),
    .io_input_mat_2(Calc6x6_1_io_input_mat_2),
    .io_input_mat_3(Calc6x6_1_io_input_mat_3),
    .io_input_mat_4(Calc6x6_1_io_input_mat_4),
    .io_input_mat_5(Calc6x6_1_io_input_mat_5),
    .io_input_mat_6(Calc6x6_1_io_input_mat_6),
    .io_input_mat_7(Calc6x6_1_io_input_mat_7),
    .io_input_mat_8(Calc6x6_1_io_input_mat_8),
    .io_input_mat_9(Calc6x6_1_io_input_mat_9),
    .io_input_mat_10(Calc6x6_1_io_input_mat_10),
    .io_input_mat_11(Calc6x6_1_io_input_mat_11),
    .io_input_mat_12(Calc6x6_1_io_input_mat_12),
    .io_input_mat_13(Calc6x6_1_io_input_mat_13),
    .io_input_mat_14(Calc6x6_1_io_input_mat_14),
    .io_input_mat_15(Calc6x6_1_io_input_mat_15),
    .io_input_mat_16(Calc6x6_1_io_input_mat_16),
    .io_input_mat_17(Calc6x6_1_io_input_mat_17),
    .io_input_mat_18(Calc6x6_1_io_input_mat_18),
    .io_input_mat_19(Calc6x6_1_io_input_mat_19),
    .io_input_mat_20(Calc6x6_1_io_input_mat_20),
    .io_input_mat_21(Calc6x6_1_io_input_mat_21),
    .io_input_mat_22(Calc6x6_1_io_input_mat_22),
    .io_input_mat_23(Calc6x6_1_io_input_mat_23),
    .io_input_mat_24(Calc6x6_1_io_input_mat_24),
    .io_input_mat_25(Calc6x6_1_io_input_mat_25),
    .io_input_mat_26(Calc6x6_1_io_input_mat_26),
    .io_input_mat_27(Calc6x6_1_io_input_mat_27),
    .io_input_mat_28(Calc6x6_1_io_input_mat_28),
    .io_input_mat_29(Calc6x6_1_io_input_mat_29),
    .io_input_mat_30(Calc6x6_1_io_input_mat_30),
    .io_input_mat_31(Calc6x6_1_io_input_mat_31),
    .io_input_mat_32(Calc6x6_1_io_input_mat_32),
    .io_input_mat_33(Calc6x6_1_io_input_mat_33),
    .io_input_mat_34(Calc6x6_1_io_input_mat_34),
    .io_input_mat_35(Calc6x6_1_io_input_mat_35),
    .io_flag(Calc6x6_1_io_flag),
    .io_weight_real_0(Calc6x6_1_io_weight_real_0),
    .io_weight_real_1(Calc6x6_1_io_weight_real_1),
    .io_weight_real_2(Calc6x6_1_io_weight_real_2),
    .io_weight_real_3(Calc6x6_1_io_weight_real_3),
    .io_weight_real_4(Calc6x6_1_io_weight_real_4),
    .io_weight_real_5(Calc6x6_1_io_weight_real_5),
    .io_weight_real_6(Calc6x6_1_io_weight_real_6),
    .io_weight_real_7(Calc6x6_1_io_weight_real_7),
    .io_weight_real_8(Calc6x6_1_io_weight_real_8),
    .io_weight_real_9(Calc6x6_1_io_weight_real_9),
    .io_weight_real_10(Calc6x6_1_io_weight_real_10),
    .io_weight_real_11(Calc6x6_1_io_weight_real_11),
    .io_weight_real_12(Calc6x6_1_io_weight_real_12),
    .io_weight_real_13(Calc6x6_1_io_weight_real_13),
    .io_weight_real_14(Calc6x6_1_io_weight_real_14),
    .io_weight_real_15(Calc6x6_1_io_weight_real_15),
    .io_weight_comp1_0(Calc6x6_1_io_weight_comp1_0),
    .io_weight_comp1_1(Calc6x6_1_io_weight_comp1_1),
    .io_weight_comp1_2(Calc6x6_1_io_weight_comp1_2),
    .io_weight_comp1_3(Calc6x6_1_io_weight_comp1_3),
    .io_weight_comp1_4(Calc6x6_1_io_weight_comp1_4),
    .io_weight_comp1_5(Calc6x6_1_io_weight_comp1_5),
    .io_weight_comp1_6(Calc6x6_1_io_weight_comp1_6),
    .io_weight_comp1_7(Calc6x6_1_io_weight_comp1_7),
    .io_weight_comp1_8(Calc6x6_1_io_weight_comp1_8),
    .io_weight_comp1_9(Calc6x6_1_io_weight_comp1_9),
    .io_weight_comp2_0(Calc6x6_1_io_weight_comp2_0),
    .io_weight_comp2_1(Calc6x6_1_io_weight_comp2_1),
    .io_weight_comp2_2(Calc6x6_1_io_weight_comp2_2),
    .io_weight_comp2_3(Calc6x6_1_io_weight_comp2_3),
    .io_weight_comp2_4(Calc6x6_1_io_weight_comp2_4),
    .io_weight_comp2_5(Calc6x6_1_io_weight_comp2_5),
    .io_weight_comp2_6(Calc6x6_1_io_weight_comp2_6),
    .io_weight_comp2_7(Calc6x6_1_io_weight_comp2_7),
    .io_weight_comp2_8(Calc6x6_1_io_weight_comp2_8),
    .io_weight_comp2_9(Calc6x6_1_io_weight_comp2_9),
    .io_weight_comp3_0(Calc6x6_1_io_weight_comp3_0),
    .io_weight_comp3_1(Calc6x6_1_io_weight_comp3_1),
    .io_weight_comp3_2(Calc6x6_1_io_weight_comp3_2),
    .io_weight_comp3_3(Calc6x6_1_io_weight_comp3_3),
    .io_weight_comp3_4(Calc6x6_1_io_weight_comp3_4),
    .io_weight_comp3_5(Calc6x6_1_io_weight_comp3_5),
    .io_weight_comp3_6(Calc6x6_1_io_weight_comp3_6),
    .io_weight_comp3_7(Calc6x6_1_io_weight_comp3_7),
    .io_weight_comp3_8(Calc6x6_1_io_weight_comp3_8),
    .io_weight_comp3_9(Calc6x6_1_io_weight_comp3_9),
    .io_output_mat_0(Calc6x6_1_io_output_mat_0),
    .io_output_mat_1(Calc6x6_1_io_output_mat_1),
    .io_output_mat_2(Calc6x6_1_io_output_mat_2),
    .io_output_mat_3(Calc6x6_1_io_output_mat_3),
    .io_output_mat_4(Calc6x6_1_io_output_mat_4),
    .io_output_mat_5(Calc6x6_1_io_output_mat_5),
    .io_output_mat_6(Calc6x6_1_io_output_mat_6),
    .io_output_mat_7(Calc6x6_1_io_output_mat_7),
    .io_output_mat_8(Calc6x6_1_io_output_mat_8),
    .io_output_mat_9(Calc6x6_1_io_output_mat_9),
    .io_output_mat_10(Calc6x6_1_io_output_mat_10),
    .io_output_mat_11(Calc6x6_1_io_output_mat_11),
    .io_output_mat_12(Calc6x6_1_io_output_mat_12),
    .io_output_mat_13(Calc6x6_1_io_output_mat_13),
    .io_output_mat_14(Calc6x6_1_io_output_mat_14),
    .io_output_mat_15(Calc6x6_1_io_output_mat_15),
    .io_valid_in(Calc6x6_1_io_valid_in),
    .io_valid_out(Calc6x6_1_io_valid_out)
  );
  Calc6x6 Calc6x6_2 ( // @[calc8x8.scala 59:39]
    .clock(Calc6x6_2_clock),
    .reset(Calc6x6_2_reset),
    .io_input_mat_0(Calc6x6_2_io_input_mat_0),
    .io_input_mat_1(Calc6x6_2_io_input_mat_1),
    .io_input_mat_2(Calc6x6_2_io_input_mat_2),
    .io_input_mat_3(Calc6x6_2_io_input_mat_3),
    .io_input_mat_4(Calc6x6_2_io_input_mat_4),
    .io_input_mat_5(Calc6x6_2_io_input_mat_5),
    .io_input_mat_6(Calc6x6_2_io_input_mat_6),
    .io_input_mat_7(Calc6x6_2_io_input_mat_7),
    .io_input_mat_8(Calc6x6_2_io_input_mat_8),
    .io_input_mat_9(Calc6x6_2_io_input_mat_9),
    .io_input_mat_10(Calc6x6_2_io_input_mat_10),
    .io_input_mat_11(Calc6x6_2_io_input_mat_11),
    .io_input_mat_12(Calc6x6_2_io_input_mat_12),
    .io_input_mat_13(Calc6x6_2_io_input_mat_13),
    .io_input_mat_14(Calc6x6_2_io_input_mat_14),
    .io_input_mat_15(Calc6x6_2_io_input_mat_15),
    .io_input_mat_16(Calc6x6_2_io_input_mat_16),
    .io_input_mat_17(Calc6x6_2_io_input_mat_17),
    .io_input_mat_18(Calc6x6_2_io_input_mat_18),
    .io_input_mat_19(Calc6x6_2_io_input_mat_19),
    .io_input_mat_20(Calc6x6_2_io_input_mat_20),
    .io_input_mat_21(Calc6x6_2_io_input_mat_21),
    .io_input_mat_22(Calc6x6_2_io_input_mat_22),
    .io_input_mat_23(Calc6x6_2_io_input_mat_23),
    .io_input_mat_24(Calc6x6_2_io_input_mat_24),
    .io_input_mat_25(Calc6x6_2_io_input_mat_25),
    .io_input_mat_26(Calc6x6_2_io_input_mat_26),
    .io_input_mat_27(Calc6x6_2_io_input_mat_27),
    .io_input_mat_28(Calc6x6_2_io_input_mat_28),
    .io_input_mat_29(Calc6x6_2_io_input_mat_29),
    .io_input_mat_30(Calc6x6_2_io_input_mat_30),
    .io_input_mat_31(Calc6x6_2_io_input_mat_31),
    .io_input_mat_32(Calc6x6_2_io_input_mat_32),
    .io_input_mat_33(Calc6x6_2_io_input_mat_33),
    .io_input_mat_34(Calc6x6_2_io_input_mat_34),
    .io_input_mat_35(Calc6x6_2_io_input_mat_35),
    .io_flag(Calc6x6_2_io_flag),
    .io_weight_real_0(Calc6x6_2_io_weight_real_0),
    .io_weight_real_1(Calc6x6_2_io_weight_real_1),
    .io_weight_real_2(Calc6x6_2_io_weight_real_2),
    .io_weight_real_3(Calc6x6_2_io_weight_real_3),
    .io_weight_real_4(Calc6x6_2_io_weight_real_4),
    .io_weight_real_5(Calc6x6_2_io_weight_real_5),
    .io_weight_real_6(Calc6x6_2_io_weight_real_6),
    .io_weight_real_7(Calc6x6_2_io_weight_real_7),
    .io_weight_real_8(Calc6x6_2_io_weight_real_8),
    .io_weight_real_9(Calc6x6_2_io_weight_real_9),
    .io_weight_real_10(Calc6x6_2_io_weight_real_10),
    .io_weight_real_11(Calc6x6_2_io_weight_real_11),
    .io_weight_real_12(Calc6x6_2_io_weight_real_12),
    .io_weight_real_13(Calc6x6_2_io_weight_real_13),
    .io_weight_real_14(Calc6x6_2_io_weight_real_14),
    .io_weight_real_15(Calc6x6_2_io_weight_real_15),
    .io_weight_comp1_0(Calc6x6_2_io_weight_comp1_0),
    .io_weight_comp1_1(Calc6x6_2_io_weight_comp1_1),
    .io_weight_comp1_2(Calc6x6_2_io_weight_comp1_2),
    .io_weight_comp1_3(Calc6x6_2_io_weight_comp1_3),
    .io_weight_comp1_4(Calc6x6_2_io_weight_comp1_4),
    .io_weight_comp1_5(Calc6x6_2_io_weight_comp1_5),
    .io_weight_comp1_6(Calc6x6_2_io_weight_comp1_6),
    .io_weight_comp1_7(Calc6x6_2_io_weight_comp1_7),
    .io_weight_comp1_8(Calc6x6_2_io_weight_comp1_8),
    .io_weight_comp1_9(Calc6x6_2_io_weight_comp1_9),
    .io_weight_comp2_0(Calc6x6_2_io_weight_comp2_0),
    .io_weight_comp2_1(Calc6x6_2_io_weight_comp2_1),
    .io_weight_comp2_2(Calc6x6_2_io_weight_comp2_2),
    .io_weight_comp2_3(Calc6x6_2_io_weight_comp2_3),
    .io_weight_comp2_4(Calc6x6_2_io_weight_comp2_4),
    .io_weight_comp2_5(Calc6x6_2_io_weight_comp2_5),
    .io_weight_comp2_6(Calc6x6_2_io_weight_comp2_6),
    .io_weight_comp2_7(Calc6x6_2_io_weight_comp2_7),
    .io_weight_comp2_8(Calc6x6_2_io_weight_comp2_8),
    .io_weight_comp2_9(Calc6x6_2_io_weight_comp2_9),
    .io_weight_comp3_0(Calc6x6_2_io_weight_comp3_0),
    .io_weight_comp3_1(Calc6x6_2_io_weight_comp3_1),
    .io_weight_comp3_2(Calc6x6_2_io_weight_comp3_2),
    .io_weight_comp3_3(Calc6x6_2_io_weight_comp3_3),
    .io_weight_comp3_4(Calc6x6_2_io_weight_comp3_4),
    .io_weight_comp3_5(Calc6x6_2_io_weight_comp3_5),
    .io_weight_comp3_6(Calc6x6_2_io_weight_comp3_6),
    .io_weight_comp3_7(Calc6x6_2_io_weight_comp3_7),
    .io_weight_comp3_8(Calc6x6_2_io_weight_comp3_8),
    .io_weight_comp3_9(Calc6x6_2_io_weight_comp3_9),
    .io_output_mat_0(Calc6x6_2_io_output_mat_0),
    .io_output_mat_1(Calc6x6_2_io_output_mat_1),
    .io_output_mat_2(Calc6x6_2_io_output_mat_2),
    .io_output_mat_3(Calc6x6_2_io_output_mat_3),
    .io_output_mat_4(Calc6x6_2_io_output_mat_4),
    .io_output_mat_5(Calc6x6_2_io_output_mat_5),
    .io_output_mat_6(Calc6x6_2_io_output_mat_6),
    .io_output_mat_7(Calc6x6_2_io_output_mat_7),
    .io_output_mat_8(Calc6x6_2_io_output_mat_8),
    .io_output_mat_9(Calc6x6_2_io_output_mat_9),
    .io_output_mat_10(Calc6x6_2_io_output_mat_10),
    .io_output_mat_11(Calc6x6_2_io_output_mat_11),
    .io_output_mat_12(Calc6x6_2_io_output_mat_12),
    .io_output_mat_13(Calc6x6_2_io_output_mat_13),
    .io_output_mat_14(Calc6x6_2_io_output_mat_14),
    .io_output_mat_15(Calc6x6_2_io_output_mat_15),
    .io_valid_in(Calc6x6_2_io_valid_in),
    .io_valid_out(Calc6x6_2_io_valid_out)
  );
  Calc6x6 Calc6x6_3 ( // @[calc8x8.scala 59:39]
    .clock(Calc6x6_3_clock),
    .reset(Calc6x6_3_reset),
    .io_input_mat_0(Calc6x6_3_io_input_mat_0),
    .io_input_mat_1(Calc6x6_3_io_input_mat_1),
    .io_input_mat_2(Calc6x6_3_io_input_mat_2),
    .io_input_mat_3(Calc6x6_3_io_input_mat_3),
    .io_input_mat_4(Calc6x6_3_io_input_mat_4),
    .io_input_mat_5(Calc6x6_3_io_input_mat_5),
    .io_input_mat_6(Calc6x6_3_io_input_mat_6),
    .io_input_mat_7(Calc6x6_3_io_input_mat_7),
    .io_input_mat_8(Calc6x6_3_io_input_mat_8),
    .io_input_mat_9(Calc6x6_3_io_input_mat_9),
    .io_input_mat_10(Calc6x6_3_io_input_mat_10),
    .io_input_mat_11(Calc6x6_3_io_input_mat_11),
    .io_input_mat_12(Calc6x6_3_io_input_mat_12),
    .io_input_mat_13(Calc6x6_3_io_input_mat_13),
    .io_input_mat_14(Calc6x6_3_io_input_mat_14),
    .io_input_mat_15(Calc6x6_3_io_input_mat_15),
    .io_input_mat_16(Calc6x6_3_io_input_mat_16),
    .io_input_mat_17(Calc6x6_3_io_input_mat_17),
    .io_input_mat_18(Calc6x6_3_io_input_mat_18),
    .io_input_mat_19(Calc6x6_3_io_input_mat_19),
    .io_input_mat_20(Calc6x6_3_io_input_mat_20),
    .io_input_mat_21(Calc6x6_3_io_input_mat_21),
    .io_input_mat_22(Calc6x6_3_io_input_mat_22),
    .io_input_mat_23(Calc6x6_3_io_input_mat_23),
    .io_input_mat_24(Calc6x6_3_io_input_mat_24),
    .io_input_mat_25(Calc6x6_3_io_input_mat_25),
    .io_input_mat_26(Calc6x6_3_io_input_mat_26),
    .io_input_mat_27(Calc6x6_3_io_input_mat_27),
    .io_input_mat_28(Calc6x6_3_io_input_mat_28),
    .io_input_mat_29(Calc6x6_3_io_input_mat_29),
    .io_input_mat_30(Calc6x6_3_io_input_mat_30),
    .io_input_mat_31(Calc6x6_3_io_input_mat_31),
    .io_input_mat_32(Calc6x6_3_io_input_mat_32),
    .io_input_mat_33(Calc6x6_3_io_input_mat_33),
    .io_input_mat_34(Calc6x6_3_io_input_mat_34),
    .io_input_mat_35(Calc6x6_3_io_input_mat_35),
    .io_flag(Calc6x6_3_io_flag),
    .io_weight_real_0(Calc6x6_3_io_weight_real_0),
    .io_weight_real_1(Calc6x6_3_io_weight_real_1),
    .io_weight_real_2(Calc6x6_3_io_weight_real_2),
    .io_weight_real_3(Calc6x6_3_io_weight_real_3),
    .io_weight_real_4(Calc6x6_3_io_weight_real_4),
    .io_weight_real_5(Calc6x6_3_io_weight_real_5),
    .io_weight_real_6(Calc6x6_3_io_weight_real_6),
    .io_weight_real_7(Calc6x6_3_io_weight_real_7),
    .io_weight_real_8(Calc6x6_3_io_weight_real_8),
    .io_weight_real_9(Calc6x6_3_io_weight_real_9),
    .io_weight_real_10(Calc6x6_3_io_weight_real_10),
    .io_weight_real_11(Calc6x6_3_io_weight_real_11),
    .io_weight_real_12(Calc6x6_3_io_weight_real_12),
    .io_weight_real_13(Calc6x6_3_io_weight_real_13),
    .io_weight_real_14(Calc6x6_3_io_weight_real_14),
    .io_weight_real_15(Calc6x6_3_io_weight_real_15),
    .io_weight_comp1_0(Calc6x6_3_io_weight_comp1_0),
    .io_weight_comp1_1(Calc6x6_3_io_weight_comp1_1),
    .io_weight_comp1_2(Calc6x6_3_io_weight_comp1_2),
    .io_weight_comp1_3(Calc6x6_3_io_weight_comp1_3),
    .io_weight_comp1_4(Calc6x6_3_io_weight_comp1_4),
    .io_weight_comp1_5(Calc6x6_3_io_weight_comp1_5),
    .io_weight_comp1_6(Calc6x6_3_io_weight_comp1_6),
    .io_weight_comp1_7(Calc6x6_3_io_weight_comp1_7),
    .io_weight_comp1_8(Calc6x6_3_io_weight_comp1_8),
    .io_weight_comp1_9(Calc6x6_3_io_weight_comp1_9),
    .io_weight_comp2_0(Calc6x6_3_io_weight_comp2_0),
    .io_weight_comp2_1(Calc6x6_3_io_weight_comp2_1),
    .io_weight_comp2_2(Calc6x6_3_io_weight_comp2_2),
    .io_weight_comp2_3(Calc6x6_3_io_weight_comp2_3),
    .io_weight_comp2_4(Calc6x6_3_io_weight_comp2_4),
    .io_weight_comp2_5(Calc6x6_3_io_weight_comp2_5),
    .io_weight_comp2_6(Calc6x6_3_io_weight_comp2_6),
    .io_weight_comp2_7(Calc6x6_3_io_weight_comp2_7),
    .io_weight_comp2_8(Calc6x6_3_io_weight_comp2_8),
    .io_weight_comp2_9(Calc6x6_3_io_weight_comp2_9),
    .io_weight_comp3_0(Calc6x6_3_io_weight_comp3_0),
    .io_weight_comp3_1(Calc6x6_3_io_weight_comp3_1),
    .io_weight_comp3_2(Calc6x6_3_io_weight_comp3_2),
    .io_weight_comp3_3(Calc6x6_3_io_weight_comp3_3),
    .io_weight_comp3_4(Calc6x6_3_io_weight_comp3_4),
    .io_weight_comp3_5(Calc6x6_3_io_weight_comp3_5),
    .io_weight_comp3_6(Calc6x6_3_io_weight_comp3_6),
    .io_weight_comp3_7(Calc6x6_3_io_weight_comp3_7),
    .io_weight_comp3_8(Calc6x6_3_io_weight_comp3_8),
    .io_weight_comp3_9(Calc6x6_3_io_weight_comp3_9),
    .io_output_mat_0(Calc6x6_3_io_output_mat_0),
    .io_output_mat_1(Calc6x6_3_io_output_mat_1),
    .io_output_mat_2(Calc6x6_3_io_output_mat_2),
    .io_output_mat_3(Calc6x6_3_io_output_mat_3),
    .io_output_mat_4(Calc6x6_3_io_output_mat_4),
    .io_output_mat_5(Calc6x6_3_io_output_mat_5),
    .io_output_mat_6(Calc6x6_3_io_output_mat_6),
    .io_output_mat_7(Calc6x6_3_io_output_mat_7),
    .io_output_mat_8(Calc6x6_3_io_output_mat_8),
    .io_output_mat_9(Calc6x6_3_io_output_mat_9),
    .io_output_mat_10(Calc6x6_3_io_output_mat_10),
    .io_output_mat_11(Calc6x6_3_io_output_mat_11),
    .io_output_mat_12(Calc6x6_3_io_output_mat_12),
    .io_output_mat_13(Calc6x6_3_io_output_mat_13),
    .io_output_mat_14(Calc6x6_3_io_output_mat_14),
    .io_output_mat_15(Calc6x6_3_io_output_mat_15),
    .io_valid_in(Calc6x6_3_io_valid_in),
    .io_valid_out(Calc6x6_3_io_valid_out)
  );
  assign io_output_mat_0 = _T_2 ? $signed(A_0_output_mat_0) : $signed(_GEN_611); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_1 = _T_2 ? $signed(A_0_output_mat_1) : $signed(_GEN_612); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_2 = _T_2 ? $signed(A_0_output_mat_2) : $signed(_GEN_613); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_3 = _T_2 ? $signed(A_0_output_mat_3) : $signed(_GEN_614); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_4 = _T_2 ? $signed(A_1_output_mat_0) : $signed(_GEN_615); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_5 = _T_2 ? $signed(A_1_output_mat_1) : $signed(_GEN_616); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_6 = _T_2 ? $signed(A_1_output_mat_2) : $signed(_GEN_617); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_7 = _T_2 ? $signed(A_1_output_mat_3) : $signed(_GEN_618); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_8 = _T_2 ? $signed(A_0_output_mat_4) : $signed(_GEN_619); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_9 = _T_2 ? $signed(A_0_output_mat_5) : $signed(_GEN_620); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_10 = _T_2 ? $signed(A_0_output_mat_6) : $signed(_GEN_621); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_11 = _T_2 ? $signed(A_0_output_mat_7) : $signed(_GEN_622); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_12 = _T_2 ? $signed(A_1_output_mat_4) : $signed(_GEN_623); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_13 = _T_2 ? $signed(A_1_output_mat_5) : $signed(_GEN_624); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_14 = _T_2 ? $signed(A_1_output_mat_6) : $signed(_GEN_625); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_15 = _T_2 ? $signed(A_1_output_mat_7) : $signed(_GEN_626); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_16 = _T_2 ? $signed(A_0_output_mat_8) : $signed(_GEN_627); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_17 = _T_2 ? $signed(A_0_output_mat_9) : $signed(_GEN_628); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_18 = _T_2 ? $signed(A_0_output_mat_10) : $signed(_GEN_629); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_19 = _T_2 ? $signed(A_0_output_mat_11) : $signed(_GEN_630); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_20 = _T_2 ? $signed(A_1_output_mat_8) : $signed(_GEN_631); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_21 = _T_2 ? $signed(A_1_output_mat_9) : $signed(_GEN_632); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_22 = _T_2 ? $signed(A_1_output_mat_10) : $signed(_GEN_633); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_23 = _T_2 ? $signed(A_1_output_mat_11) : $signed(_GEN_634); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_24 = _T_2 ? $signed(A_0_output_mat_12) : $signed(_GEN_635); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_25 = _T_2 ? $signed(A_0_output_mat_13) : $signed(_GEN_636); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_26 = _T_2 ? $signed(A_0_output_mat_14) : $signed(_GEN_637); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_27 = _T_2 ? $signed(A_0_output_mat_15) : $signed(_GEN_638); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_28 = _T_2 ? $signed(A_1_output_mat_12) : $signed(_GEN_639); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_29 = _T_2 ? $signed(A_1_output_mat_13) : $signed(_GEN_640); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_30 = _T_2 ? $signed(A_1_output_mat_14) : $signed(_GEN_641); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_31 = _T_2 ? $signed(A_1_output_mat_15) : $signed(_GEN_642); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_32 = _T_2 ? $signed(A_2_output_mat_0) : $signed(_GEN_643); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_33 = _T_2 ? $signed(A_2_output_mat_1) : $signed(_GEN_644); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_34 = _T_2 ? $signed(A_2_output_mat_2) : $signed(_GEN_645); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_35 = _T_2 ? $signed(A_2_output_mat_3) : $signed(_GEN_646); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_36 = _T_2 ? $signed(A_3_output_mat_0) : $signed(_GEN_647); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_37 = _T_2 ? $signed(A_3_output_mat_1) : $signed(_GEN_648); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_38 = _T_2 ? $signed(A_3_output_mat_2) : $signed(_GEN_649); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_39 = _T_2 ? $signed(A_3_output_mat_3) : $signed(_GEN_650); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_40 = _T_2 ? $signed(A_2_output_mat_4) : $signed(_GEN_651); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_41 = _T_2 ? $signed(A_2_output_mat_5) : $signed(_GEN_652); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_42 = _T_2 ? $signed(A_2_output_mat_6) : $signed(_GEN_653); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_43 = _T_2 ? $signed(A_2_output_mat_7) : $signed(_GEN_654); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_44 = _T_2 ? $signed(A_3_output_mat_4) : $signed(_GEN_655); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_45 = _T_2 ? $signed(A_3_output_mat_5) : $signed(_GEN_656); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_46 = _T_2 ? $signed(A_3_output_mat_6) : $signed(_GEN_657); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_47 = _T_2 ? $signed(A_3_output_mat_7) : $signed(_GEN_658); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_48 = _T_2 ? $signed(A_2_output_mat_8) : $signed(_GEN_659); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_49 = _T_2 ? $signed(A_2_output_mat_9) : $signed(_GEN_660); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_50 = _T_2 ? $signed(A_2_output_mat_10) : $signed(_GEN_661); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_51 = _T_2 ? $signed(A_2_output_mat_11) : $signed(_GEN_662); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_52 = _T_2 ? $signed(A_3_output_mat_8) : $signed(_GEN_663); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_53 = _T_2 ? $signed(A_3_output_mat_9) : $signed(_GEN_664); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_54 = _T_2 ? $signed(A_3_output_mat_10) : $signed(_GEN_665); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_55 = _T_2 ? $signed(A_3_output_mat_11) : $signed(_GEN_666); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_56 = _T_2 ? $signed(A_2_output_mat_12) : $signed(_GEN_667); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_57 = _T_2 ? $signed(A_2_output_mat_13) : $signed(_GEN_668); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_58 = _T_2 ? $signed(A_2_output_mat_14) : $signed(_GEN_669); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_59 = _T_2 ? $signed(A_2_output_mat_15) : $signed(_GEN_670); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_60 = _T_2 ? $signed(A_3_output_mat_12) : $signed(_GEN_671); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_61 = _T_2 ? $signed(A_3_output_mat_13) : $signed(_GEN_672); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_62 = _T_2 ? $signed(A_3_output_mat_14) : $signed(_GEN_673); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_output_mat_63 = _T_2 ? $signed(A_3_output_mat_15) : $signed(_GEN_674); // @[Conditional.scala 40:58 calc8x8.scala 146:23]
  assign io_valid_out = _T_2 ? A_0_valid_out : _GEN_675; // @[Conditional.scala 40:58 calc8x8.scala 147:26]
  assign Calc6x6_clock = clock;
  assign Calc6x6_reset = reset;
  assign Calc6x6_io_input_mat_0 = _T_2 ? $signed(io_input_mat_0) : $signed(_GEN_398); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_1 = _T_2 ? $signed(io_input_mat_1) : $signed(_GEN_399); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_2 = _T_2 ? $signed(io_input_mat_2) : $signed(_GEN_400); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_3 = _T_2 ? $signed(io_input_mat_3) : $signed(_GEN_401); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_4 = _T_2 ? $signed(16'sh0) : $signed(_GEN_402); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_5 = _T_2 ? $signed(16'sh0) : $signed(_GEN_403); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_6 = _T_2 ? $signed(io_input_mat_8) : $signed(_GEN_404); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_7 = _T_2 ? $signed(io_input_mat_9) : $signed(_GEN_405); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_8 = _T_2 ? $signed(io_input_mat_10) : $signed(_GEN_406); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_9 = _T_2 ? $signed(io_input_mat_11) : $signed(_GEN_407); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_10 = _T_2 ? $signed(16'sh0) : $signed(_GEN_408); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_11 = _T_2 ? $signed(16'sh0) : $signed(_GEN_409); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_12 = _T_2 ? $signed(io_input_mat_16) : $signed(_GEN_410); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_13 = _T_2 ? $signed(io_input_mat_17) : $signed(_GEN_411); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_14 = _T_2 ? $signed(io_input_mat_18) : $signed(_GEN_412); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_15 = _T_2 ? $signed(io_input_mat_19) : $signed(_GEN_413); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_16 = _T_2 ? $signed(16'sh0) : $signed(_GEN_414); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_17 = _T_2 ? $signed(16'sh0) : $signed(_GEN_415); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_18 = _T_2 ? $signed(io_input_mat_24) : $signed(_GEN_416); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_19 = _T_2 ? $signed(io_input_mat_25) : $signed(_GEN_417); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_20 = _T_2 ? $signed(io_input_mat_26) : $signed(_GEN_418); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_21 = _T_2 ? $signed(io_input_mat_27) : $signed(_GEN_419); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_22 = _T_2 ? $signed(16'sh0) : $signed(_GEN_420); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_23 = _T_2 ? $signed(16'sh0) : $signed(_GEN_421); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_24 = _T_2 ? $signed(16'sh0) : $signed(_GEN_422); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_25 = _T_2 ? $signed(16'sh0) : $signed(_GEN_423); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_26 = _T_2 ? $signed(16'sh0) : $signed(_GEN_424); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_27 = _T_2 ? $signed(16'sh0) : $signed(_GEN_425); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_28 = _T_2 ? $signed(16'sh0) : $signed(_GEN_426); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_29 = _T_2 ? $signed(16'sh0) : $signed(_GEN_427); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_30 = _T_2 ? $signed(16'sh0) : $signed(_GEN_428); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_31 = _T_2 ? $signed(16'sh0) : $signed(_GEN_429); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_32 = _T_2 ? $signed(16'sh0) : $signed(_GEN_430); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_33 = _T_2 ? $signed(16'sh0) : $signed(_GEN_431); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_34 = _T_2 ? $signed(16'sh0) : $signed(_GEN_432); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_input_mat_35 = _T_2 ? $signed(16'sh0) : $signed(_GEN_433); // @[Conditional.scala 40:58 calc8x8.scala 138:24]
  assign Calc6x6_io_flag = _T_2 ? 2'h0 : _GEN_558; // @[Conditional.scala 40:58 calc8x8.scala 143:27]
  assign Calc6x6_io_weight_real_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_542); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_543); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_544); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_545); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_546); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_547); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_548); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_549); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_550); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_551); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_10 = _T_2 ? $signed(18'sh0) : $signed(_GEN_552); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_11 = _T_2 ? $signed(18'sh0) : $signed(_GEN_553); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_12 = _T_2 ? $signed(18'sh0) : $signed(_GEN_554); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_13 = _T_2 ? $signed(18'sh0) : $signed(_GEN_555); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_14 = _T_2 ? $signed(18'sh0) : $signed(_GEN_556); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_real_15 = _T_2 ? $signed(18'sh0) : $signed(_GEN_557); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_696); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_697); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_698); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_699); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_700); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_701); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_702); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_703); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_704); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp1_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_705); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_686); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_687); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_688); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_689); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_690); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_691); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_692); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_693); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_694); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp2_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_695); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_676); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_677); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_678); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_679); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_680); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_681); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_682); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_683); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_684); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_weight_comp3_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_685); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_io_valid_in = _T_2 ? io_valid_in : _GEN_559; // @[Conditional.scala 40:58 calc8x8.scala 144:31]
  assign Calc6x6_1_clock = clock;
  assign Calc6x6_1_reset = reset;
  assign Calc6x6_1_io_input_mat_0 = _T_2 ? $signed(io_input_mat_3) : $signed(_GEN_434); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_1 = _T_2 ? $signed(io_input_mat_4) : $signed(_GEN_435); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_2 = _T_2 ? $signed(io_input_mat_5) : $signed(_GEN_436); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_3 = _T_2 ? $signed(io_input_mat_6) : $signed(_GEN_437); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_4 = _T_2 ? $signed(io_input_mat_7) : $signed(_GEN_438); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_5 = _T_2 ? $signed(16'sh0) : $signed(_GEN_439); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_6 = _T_2 ? $signed(io_input_mat_11) : $signed(_GEN_440); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_7 = _T_2 ? $signed(io_input_mat_12) : $signed(_GEN_441); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_8 = _T_2 ? $signed(io_input_mat_13) : $signed(_GEN_442); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_9 = _T_2 ? $signed(io_input_mat_14) : $signed(_GEN_443); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_10 = _T_2 ? $signed(io_input_mat_15) : $signed(_GEN_444); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_11 = _T_2 ? $signed(16'sh0) : $signed(_GEN_445); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_12 = _T_2 ? $signed(io_input_mat_19) : $signed(_GEN_446); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_13 = _T_2 ? $signed(io_input_mat_20) : $signed(_GEN_447); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_14 = _T_2 ? $signed(io_input_mat_21) : $signed(_GEN_448); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_15 = _T_2 ? $signed(io_input_mat_22) : $signed(_GEN_449); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_16 = _T_2 ? $signed(io_input_mat_23) : $signed(_GEN_450); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_17 = _T_2 ? $signed(16'sh0) : $signed(_GEN_451); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_18 = _T_2 ? $signed(io_input_mat_27) : $signed(_GEN_452); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_19 = _T_2 ? $signed(io_input_mat_28) : $signed(_GEN_453); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_20 = _T_2 ? $signed(io_input_mat_29) : $signed(_GEN_454); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_21 = _T_2 ? $signed(io_input_mat_30) : $signed(_GEN_455); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_22 = _T_2 ? $signed(io_input_mat_31) : $signed(_GEN_456); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_23 = _T_2 ? $signed(16'sh0) : $signed(_GEN_457); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_24 = _T_2 ? $signed(16'sh0) : $signed(_GEN_426); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_25 = _T_2 ? $signed(16'sh0) : $signed(_GEN_427); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_26 = _T_2 ? $signed(16'sh0) : $signed(_GEN_460); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_27 = _T_2 ? $signed(16'sh0) : $signed(_GEN_461); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_28 = _T_2 ? $signed(16'sh0) : $signed(_GEN_462); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_29 = _T_2 ? $signed(16'sh0) : $signed(_GEN_463); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_30 = _T_2 ? $signed(16'sh0) : $signed(_GEN_432); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_31 = _T_2 ? $signed(16'sh0) : $signed(_GEN_433); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_32 = _T_2 ? $signed(16'sh0) : $signed(_GEN_466); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_33 = _T_2 ? $signed(16'sh0) : $signed(_GEN_467); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_34 = _T_2 ? $signed(16'sh0) : $signed(_GEN_468); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_input_mat_35 = _T_2 ? $signed(16'sh0) : $signed(_GEN_469); // @[Conditional.scala 40:58 calc8x8.scala 139:24]
  assign Calc6x6_1_io_flag = _T_2 ? 2'h0 : _GEN_558; // @[Conditional.scala 40:58 calc8x8.scala 143:27]
  assign Calc6x6_1_io_weight_real_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_560); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_561); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_562); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_563); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_564); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_565); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_566); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_567); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_568); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_569); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_10 = _T_2 ? $signed(18'sh0) : $signed(_GEN_570); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_11 = _T_2 ? $signed(18'sh0) : $signed(_GEN_571); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_12 = _T_2 ? $signed(18'sh0) : $signed(_GEN_572); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_13 = _T_2 ? $signed(18'sh0) : $signed(_GEN_573); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_14 = _T_2 ? $signed(18'sh0) : $signed(_GEN_574); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_real_15 = _T_2 ? $signed(18'sh0) : $signed(_GEN_575); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_696); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_697); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_698); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_699); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_700); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_701); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_702); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_703); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_704); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp1_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_705); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_686); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_687); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_688); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_689); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_690); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_691); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_692); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_693); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_694); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp2_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_695); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_676); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_677); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_678); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_679); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_680); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_681); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_682); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_683); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_684); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_weight_comp3_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_685); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_1_io_valid_in = _T_2 ? io_valid_in : _GEN_559; // @[Conditional.scala 40:58 calc8x8.scala 144:31]
  assign Calc6x6_2_clock = clock;
  assign Calc6x6_2_reset = reset;
  assign Calc6x6_2_io_input_mat_0 = _T_2 ? $signed(io_input_mat_24) : $signed(_GEN_470); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_1 = _T_2 ? $signed(io_input_mat_25) : $signed(_GEN_471); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_2 = _T_2 ? $signed(io_input_mat_26) : $signed(_GEN_472); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_3 = _T_2 ? $signed(io_input_mat_27) : $signed(_GEN_473); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_4 = _T_2 ? $signed(16'sh0) : $signed(_GEN_426); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_5 = _T_2 ? $signed(16'sh0) : $signed(_GEN_427); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_6 = _T_2 ? $signed(io_input_mat_32) : $signed(_GEN_476); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_7 = _T_2 ? $signed(io_input_mat_33) : $signed(_GEN_477); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_8 = _T_2 ? $signed(io_input_mat_34) : $signed(_GEN_478); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_9 = _T_2 ? $signed(io_input_mat_35) : $signed(_GEN_479); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_10 = _T_2 ? $signed(16'sh0) : $signed(_GEN_432); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_11 = _T_2 ? $signed(16'sh0) : $signed(_GEN_433); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_12 = _T_2 ? $signed(io_input_mat_40) : $signed(_GEN_482); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_13 = _T_2 ? $signed(io_input_mat_41) : $signed(_GEN_483); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_14 = _T_2 ? $signed(io_input_mat_42) : $signed(_GEN_484); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_15 = _T_2 ? $signed(io_input_mat_43) : $signed(_GEN_485); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_16 = _T_2 ? $signed(16'sh0) : $signed(_GEN_486); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_17 = _T_2 ? $signed(16'sh0) : $signed(_GEN_487); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_18 = _T_2 ? $signed(io_input_mat_48) : $signed(_GEN_488); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_19 = _T_2 ? $signed(io_input_mat_49) : $signed(_GEN_489); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_20 = _T_2 ? $signed(io_input_mat_50) : $signed(_GEN_490); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_21 = _T_2 ? $signed(io_input_mat_51) : $signed(_GEN_491); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_22 = _T_2 ? $signed(16'sh0) : $signed(_GEN_492); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_23 = _T_2 ? $signed(16'sh0) : $signed(_GEN_493); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_24 = _T_2 ? $signed(io_input_mat_56) : $signed(_GEN_494); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_25 = _T_2 ? $signed(io_input_mat_57) : $signed(_GEN_495); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_26 = _T_2 ? $signed(io_input_mat_58) : $signed(_GEN_496); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_27 = _T_2 ? $signed(io_input_mat_59) : $signed(_GEN_497); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_28 = _T_2 ? $signed(16'sh0) : $signed(_GEN_498); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_29 = _T_2 ? $signed(16'sh0) : $signed(_GEN_499); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_30 = _T_2 ? $signed(16'sh0) : $signed(_GEN_500); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_31 = _T_2 ? $signed(16'sh0) : $signed(_GEN_501); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_32 = _T_2 ? $signed(16'sh0) : $signed(_GEN_502); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_33 = _T_2 ? $signed(16'sh0) : $signed(_GEN_503); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_34 = _T_2 ? $signed(16'sh0) : $signed(_GEN_504); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_input_mat_35 = _T_2 ? $signed(16'sh0) : $signed(_GEN_505); // @[Conditional.scala 40:58 calc8x8.scala 140:24]
  assign Calc6x6_2_io_flag = _T_2 ? 2'h0 : _GEN_558; // @[Conditional.scala 40:58 calc8x8.scala 143:27]
  assign Calc6x6_2_io_weight_real_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_577); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_578); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_579); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_580); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_581); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_582); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_583); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_584); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_585); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_586); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_10 = _T_2 ? $signed(18'sh0) : $signed(_GEN_587); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_11 = _T_2 ? $signed(18'sh0) : $signed(_GEN_588); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_12 = _T_2 ? $signed(18'sh0) : $signed(_GEN_589); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_13 = _T_2 ? $signed(18'sh0) : $signed(_GEN_590); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_14 = _T_2 ? $signed(18'sh0) : $signed(_GEN_591); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_real_15 = _T_2 ? $signed(18'sh0) : $signed(_GEN_592); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_696); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_697); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_698); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_699); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_700); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_701); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_702); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_703); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_704); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp1_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_705); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_686); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_687); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_688); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_689); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_690); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_691); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_692); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_693); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_694); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp2_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_695); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_676); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_677); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_678); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_679); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_680); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_681); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_682); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_683); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_684); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_weight_comp3_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_685); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_2_io_valid_in = _T_2 ? io_valid_in : _GEN_559; // @[Conditional.scala 40:58 calc8x8.scala 144:31]
  assign Calc6x6_3_clock = clock;
  assign Calc6x6_3_reset = reset;
  assign Calc6x6_3_io_input_mat_0 = _T_2 ? $signed(io_input_mat_27) : $signed(_GEN_506); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_1 = _T_2 ? $signed(io_input_mat_28) : $signed(_GEN_507); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_2 = _T_2 ? $signed(io_input_mat_29) : $signed(_GEN_508); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_3 = _T_2 ? $signed(io_input_mat_30) : $signed(_GEN_509); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_4 = _T_2 ? $signed(io_input_mat_31) : $signed(_GEN_510); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_5 = _T_2 ? $signed(16'sh0) : $signed(_GEN_463); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_6 = _T_2 ? $signed(io_input_mat_35) : $signed(_GEN_512); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_7 = _T_2 ? $signed(io_input_mat_36) : $signed(_GEN_513); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_8 = _T_2 ? $signed(io_input_mat_37) : $signed(_GEN_514); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_9 = _T_2 ? $signed(io_input_mat_38) : $signed(_GEN_515); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_10 = _T_2 ? $signed(io_input_mat_39) : $signed(_GEN_516); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_11 = _T_2 ? $signed(16'sh0) : $signed(_GEN_469); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_12 = _T_2 ? $signed(io_input_mat_43) : $signed(_GEN_518); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_13 = _T_2 ? $signed(io_input_mat_44) : $signed(_GEN_519); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_14 = _T_2 ? $signed(io_input_mat_45) : $signed(_GEN_520); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_15 = _T_2 ? $signed(io_input_mat_46) : $signed(_GEN_521); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_16 = _T_2 ? $signed(io_input_mat_47) : $signed(_GEN_522); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_17 = _T_2 ? $signed(16'sh0) : $signed(_GEN_523); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_18 = _T_2 ? $signed(io_input_mat_51) : $signed(_GEN_524); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_19 = _T_2 ? $signed(io_input_mat_52) : $signed(_GEN_525); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_20 = _T_2 ? $signed(io_input_mat_53) : $signed(_GEN_526); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_21 = _T_2 ? $signed(io_input_mat_54) : $signed(_GEN_527); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_22 = _T_2 ? $signed(io_input_mat_55) : $signed(_GEN_528); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_23 = _T_2 ? $signed(16'sh0) : $signed(_GEN_529); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_24 = _T_2 ? $signed(io_input_mat_59) : $signed(_GEN_530); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_25 = _T_2 ? $signed(io_input_mat_60) : $signed(_GEN_531); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_26 = _T_2 ? $signed(io_input_mat_61) : $signed(_GEN_532); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_27 = _T_2 ? $signed(io_input_mat_62) : $signed(_GEN_533); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_28 = _T_2 ? $signed(io_input_mat_63) : $signed(_GEN_534); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_29 = _T_2 ? $signed(16'sh0) : $signed(_GEN_535); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_30 = _T_2 ? $signed(16'sh0) : $signed(_GEN_504); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_31 = _T_2 ? $signed(16'sh0) : $signed(_GEN_505); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_32 = _T_2 ? $signed(16'sh0) : $signed(_GEN_538); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_33 = _T_2 ? $signed(16'sh0) : $signed(_GEN_539); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_34 = _T_2 ? $signed(16'sh0) : $signed(_GEN_540); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_input_mat_35 = _T_2 ? $signed(16'sh0) : $signed(_GEN_541); // @[Conditional.scala 40:58 calc8x8.scala 141:24]
  assign Calc6x6_3_io_flag = _T_2 ? 2'h0 : _GEN_558; // @[Conditional.scala 40:58 calc8x8.scala 143:27]
  assign Calc6x6_3_io_weight_real_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_594); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_595); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_596); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_597); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_598); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_599); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_600); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_601); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_602); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_603); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_10 = _T_2 ? $signed(18'sh0) : $signed(_GEN_604); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_11 = _T_2 ? $signed(18'sh0) : $signed(_GEN_605); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_12 = _T_2 ? $signed(18'sh0) : $signed(_GEN_606); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_13 = _T_2 ? $signed(18'sh0) : $signed(_GEN_607); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_14 = _T_2 ? $signed(18'sh0) : $signed(_GEN_608); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_real_15 = _T_2 ? $signed(18'sh0) : $signed(_GEN_609); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_696); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_697); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_698); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_699); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_700); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_701); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_702); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_703); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_704); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp1_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_705); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_686); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_687); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_688); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_689); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_690); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_691); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_692); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_693); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_694); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp2_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_695); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_0 = _T_2 ? $signed(18'sh0) : $signed(_GEN_676); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_1 = _T_2 ? $signed(18'sh0) : $signed(_GEN_677); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_2 = _T_2 ? $signed(18'sh0) : $signed(_GEN_678); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_3 = _T_2 ? $signed(18'sh0) : $signed(_GEN_679); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_4 = _T_2 ? $signed(18'sh0) : $signed(_GEN_680); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_5 = _T_2 ? $signed(18'sh0) : $signed(_GEN_681); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_6 = _T_2 ? $signed(18'sh0) : $signed(_GEN_682); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_7 = _T_2 ? $signed(18'sh0) : $signed(_GEN_683); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_8 = _T_2 ? $signed(18'sh0) : $signed(_GEN_684); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_weight_comp3_9 = _T_2 ? $signed(18'sh0) : $signed(_GEN_685); // @[Conditional.scala 40:58 calc8x8.scala 63:21]
  assign Calc6x6_3_io_valid_in = _T_2 ? io_valid_in : _GEN_559; // @[Conditional.scala 40:58 calc8x8.scala 144:31]
  always @(posedge clock) begin
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_0_0 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_0_0 <= {{2{io_weight_0_real_0[15]}},io_weight_0_real_0}; // @[calc8x8.scala 78:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_0_1 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_0_1 <= {{2{io_weight_0_real_1[15]}},io_weight_0_real_1}; // @[calc8x8.scala 78:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_0_2 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_0_2 <= {{2{io_weight_0_real_2[15]}},io_weight_0_real_2}; // @[calc8x8.scala 78:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_1_0 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_1_0 <= {{2{__B_1_0_T_5[15]}},__B_1_0_T_5}; // @[calc8x8.scala 79:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_1_1 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_1_1 <= {{2{__B_1_1_T_5[15]}},__B_1_1_T_5}; // @[calc8x8.scala 79:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_1_2 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_1_2 <= {{2{__B_1_2_T_5[15]}},__B_1_2_T_5}; // @[calc8x8.scala 79:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_2_0 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_2_0 <= {{2{__B_2_0_T_5[15]}},__B_2_0_T_5}; // @[calc8x8.scala 80:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_2_1 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_2_1 <= {{2{__B_2_1_T_5[15]}},__B_2_1_T_5}; // @[calc8x8.scala 80:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_2_2 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_2_2 <= {{2{__B_2_2_T_5[15]}},__B_2_2_T_5}; // @[calc8x8.scala 80:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_3_0 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_3_0 <= {{2{__B_3_0_T_2[15]}},__B_3_0_T_2}; // @[calc8x8.scala 81:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_3_1 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_3_1 <= {{2{__B_3_1_T_2[15]}},__B_3_1_T_2}; // @[calc8x8.scala 81:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_3_2 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_3_2 <= {{2{__B_3_2_T_2[15]}},__B_3_2_T_2}; // @[calc8x8.scala 81:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_5_0 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_5_0 <= {{2{io_weight_0_real_6[15]}},io_weight_0_real_6}; // @[calc8x8.scala 83:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_5_1 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_5_1 <= {{2{io_weight_0_real_7[15]}},io_weight_0_real_7}; // @[calc8x8.scala 83:18]
    end
    if (reset) begin // @[calc8x8.scala 71:21]
      _B_5_2 <= 18'sh0; // @[calc8x8.scala 71:21]
    end else begin
      _B_5_2 <= {{2{io_weight_0_real_8[15]}},io_weight_0_real_8}; // @[calc8x8.scala 83:18]
    end
    if (reset) begin // @[calc8x8.scala 72:22]
      _Bi_3_0 <= 18'sh0; // @[calc8x8.scala 72:22]
    end else begin
      _Bi_3_0 <= {{2{io_weight_0_real_3[15]}},io_weight_0_real_3}; // @[calc8x8.scala 84:19]
    end
    if (reset) begin // @[calc8x8.scala 72:22]
      _Bi_3_1 <= 18'sh0; // @[calc8x8.scala 72:22]
    end else begin
      _Bi_3_1 <= {{2{io_weight_0_real_4[15]}},io_weight_0_real_4}; // @[calc8x8.scala 84:19]
    end
    if (reset) begin // @[calc8x8.scala 72:22]
      _Bi_3_2 <= 18'sh0; // @[calc8x8.scala 72:22]
    end else begin
      _Bi_3_2 <= {{2{io_weight_0_real_5[15]}},io_weight_0_real_5}; // @[calc8x8.scala 84:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_0_0 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_0_0 <= {{1{_B_0_0[17]}},_B_0_0}; // @[calc8x8.scala 93:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_0_1 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_0_1 <= {{1{___B_0_1_T_5[17]}},___B_0_1_T_5}; // @[calc8x8.scala 94:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_0_2 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_0_2 <= {{1{___B_0_2_T_5[17]}},___B_0_2_T_5}; // @[calc8x8.scala 95:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_0_3 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_0_3 <= {{1{___B_0_3_T_5[17]}},___B_0_3_T_5}; // @[calc8x8.scala 96:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_0_5 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_0_5 <= {{1{_B_0_2[17]}},_B_0_2}; // @[calc8x8.scala 98:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_1_0 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_1_0 <= {{1{_B_1_0[17]}},_B_1_0}; // @[calc8x8.scala 93:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_1_1 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_1_1 <= {{1{___B_1_1_T_5[17]}},___B_1_1_T_5}; // @[calc8x8.scala 94:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_1_2 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_1_2 <= {{1{___B_1_2_T_5[17]}},___B_1_2_T_5}; // @[calc8x8.scala 95:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_1_3 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_1_3 <= {{1{___B_1_3_T_5[17]}},___B_1_3_T_5}; // @[calc8x8.scala 96:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_1_5 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_1_5 <= {{1{_B_1_2[17]}},_B_1_2}; // @[calc8x8.scala 98:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_2_0 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_2_0 <= {{1{_B_2_0[17]}},_B_2_0}; // @[calc8x8.scala 93:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_2_1 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_2_1 <= {{1{___B_2_1_T_5[17]}},___B_2_1_T_5}; // @[calc8x8.scala 94:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_2_2 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_2_2 <= {{1{___B_2_2_T_5[17]}},___B_2_2_T_5}; // @[calc8x8.scala 95:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_2_3 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_2_3 <= {{1{___B_2_3_T_5[17]}},___B_2_3_T_5}; // @[calc8x8.scala 96:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_2_5 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_2_5 <= {{1{_B_2_2[17]}},_B_2_2}; // @[calc8x8.scala 98:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_3_0 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_3_0 <= {{1{_B_3_0[17]}},_B_3_0}; // @[calc8x8.scala 93:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_3_1 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_3_1 <= {{1{___B_3_1_T_5[17]}},___B_3_1_T_5}; // @[calc8x8.scala 94:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_3_2 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_3_2 <= {{1{___B_3_2_T_5[17]}},___B_3_2_T_5}; // @[calc8x8.scala 95:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_3_3 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_3_3 <= {{1{___B_3_3_T_5[17]}},___B_3_3_T_5}; // @[calc8x8.scala 96:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_3_4 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_3_4 <= {{1{___B_3_4_T_5[17]}},___B_3_4_T_5}; // @[calc8x8.scala 97:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_3_5 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_3_5 <= {{1{_B_3_2[17]}},_B_3_2}; // @[calc8x8.scala 98:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_5_0 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_5_0 <= {{1{_B_5_0[17]}},_B_5_0}; // @[calc8x8.scala 93:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_5_1 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_5_1 <= {{1{___B_5_1_T_5[17]}},___B_5_1_T_5}; // @[calc8x8.scala 94:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_5_2 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_5_2 <= {{1{___B_5_2_T_5[17]}},___B_5_2_T_5}; // @[calc8x8.scala 95:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_5_3 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_5_3 <= {{1{___B_5_3_T_5[17]}},___B_5_3_T_5}; // @[calc8x8.scala 96:19]
    end
    if (reset) begin // @[calc8x8.scala 89:22]
      __B_5_5 <= 19'sh0; // @[calc8x8.scala 89:22]
    end else begin
      __B_5_5 <= {{1{_B_5_2[17]}},_B_5_2}; // @[calc8x8.scala 98:19]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_0_3 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_0_3 <= {{1{___Bi_0_3_T_5[17]}},___Bi_0_3_T_5}; // @[calc8x8.scala 102:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_1_3 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_1_3 <= {{1{___Bi_1_3_T_5[17]}},___Bi_1_3_T_5}; // @[calc8x8.scala 102:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_2_3 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_2_3 <= {{1{___Bi_2_3_T_5[17]}},___Bi_2_3_T_5}; // @[calc8x8.scala 102:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_3_0 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_3_0 <= {{1{_Bi_3_0[17]}},_Bi_3_0}; // @[calc8x8.scala 99:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_3_1 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_3_1 <= {{1{___Bi_3_1_T_5[17]}},___Bi_3_1_T_5}; // @[calc8x8.scala 100:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_3_2 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_3_2 <= {{1{___Bi_3_2_T_5[17]}},___Bi_3_2_T_5}; // @[calc8x8.scala 101:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_3_3 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_3_3 <= {{1{___Bi_3_3_T_5[17]}},___Bi_3_3_T_5}; // @[calc8x8.scala 102:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_3_4 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_3_4 <= {{1{___Bi_3_4_T_5[17]}},___Bi_3_4_T_5}; // @[calc8x8.scala 103:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_3_5 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_3_5 <= {{1{_Bi_3_2[17]}},_Bi_3_2}; // @[calc8x8.scala 104:20]
    end
    if (reset) begin // @[calc8x8.scala 90:23]
      __Bi_5_3 <= 19'sh0; // @[calc8x8.scala 90:23]
    end else begin
      __Bi_5_3 <= {{1{___Bi_5_3_T_5[17]}},___Bi_5_3_T_5}; // @[calc8x8.scala 102:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _B_0_0 = _RAND_0[17:0];
  _RAND_1 = {1{`RANDOM}};
  _B_0_1 = _RAND_1[17:0];
  _RAND_2 = {1{`RANDOM}};
  _B_0_2 = _RAND_2[17:0];
  _RAND_3 = {1{`RANDOM}};
  _B_1_0 = _RAND_3[17:0];
  _RAND_4 = {1{`RANDOM}};
  _B_1_1 = _RAND_4[17:0];
  _RAND_5 = {1{`RANDOM}};
  _B_1_2 = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  _B_2_0 = _RAND_6[17:0];
  _RAND_7 = {1{`RANDOM}};
  _B_2_1 = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  _B_2_2 = _RAND_8[17:0];
  _RAND_9 = {1{`RANDOM}};
  _B_3_0 = _RAND_9[17:0];
  _RAND_10 = {1{`RANDOM}};
  _B_3_1 = _RAND_10[17:0];
  _RAND_11 = {1{`RANDOM}};
  _B_3_2 = _RAND_11[17:0];
  _RAND_12 = {1{`RANDOM}};
  _B_5_0 = _RAND_12[17:0];
  _RAND_13 = {1{`RANDOM}};
  _B_5_1 = _RAND_13[17:0];
  _RAND_14 = {1{`RANDOM}};
  _B_5_2 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  _Bi_3_0 = _RAND_15[17:0];
  _RAND_16 = {1{`RANDOM}};
  _Bi_3_1 = _RAND_16[17:0];
  _RAND_17 = {1{`RANDOM}};
  _Bi_3_2 = _RAND_17[17:0];
  _RAND_18 = {1{`RANDOM}};
  __B_0_0 = _RAND_18[18:0];
  _RAND_19 = {1{`RANDOM}};
  __B_0_1 = _RAND_19[18:0];
  _RAND_20 = {1{`RANDOM}};
  __B_0_2 = _RAND_20[18:0];
  _RAND_21 = {1{`RANDOM}};
  __B_0_3 = _RAND_21[18:0];
  _RAND_22 = {1{`RANDOM}};
  __B_0_5 = _RAND_22[18:0];
  _RAND_23 = {1{`RANDOM}};
  __B_1_0 = _RAND_23[18:0];
  _RAND_24 = {1{`RANDOM}};
  __B_1_1 = _RAND_24[18:0];
  _RAND_25 = {1{`RANDOM}};
  __B_1_2 = _RAND_25[18:0];
  _RAND_26 = {1{`RANDOM}};
  __B_1_3 = _RAND_26[18:0];
  _RAND_27 = {1{`RANDOM}};
  __B_1_5 = _RAND_27[18:0];
  _RAND_28 = {1{`RANDOM}};
  __B_2_0 = _RAND_28[18:0];
  _RAND_29 = {1{`RANDOM}};
  __B_2_1 = _RAND_29[18:0];
  _RAND_30 = {1{`RANDOM}};
  __B_2_2 = _RAND_30[18:0];
  _RAND_31 = {1{`RANDOM}};
  __B_2_3 = _RAND_31[18:0];
  _RAND_32 = {1{`RANDOM}};
  __B_2_5 = _RAND_32[18:0];
  _RAND_33 = {1{`RANDOM}};
  __B_3_0 = _RAND_33[18:0];
  _RAND_34 = {1{`RANDOM}};
  __B_3_1 = _RAND_34[18:0];
  _RAND_35 = {1{`RANDOM}};
  __B_3_2 = _RAND_35[18:0];
  _RAND_36 = {1{`RANDOM}};
  __B_3_3 = _RAND_36[18:0];
  _RAND_37 = {1{`RANDOM}};
  __B_3_4 = _RAND_37[18:0];
  _RAND_38 = {1{`RANDOM}};
  __B_3_5 = _RAND_38[18:0];
  _RAND_39 = {1{`RANDOM}};
  __B_5_0 = _RAND_39[18:0];
  _RAND_40 = {1{`RANDOM}};
  __B_5_1 = _RAND_40[18:0];
  _RAND_41 = {1{`RANDOM}};
  __B_5_2 = _RAND_41[18:0];
  _RAND_42 = {1{`RANDOM}};
  __B_5_3 = _RAND_42[18:0];
  _RAND_43 = {1{`RANDOM}};
  __B_5_5 = _RAND_43[18:0];
  _RAND_44 = {1{`RANDOM}};
  __Bi_0_3 = _RAND_44[18:0];
  _RAND_45 = {1{`RANDOM}};
  __Bi_1_3 = _RAND_45[18:0];
  _RAND_46 = {1{`RANDOM}};
  __Bi_2_3 = _RAND_46[18:0];
  _RAND_47 = {1{`RANDOM}};
  __Bi_3_0 = _RAND_47[18:0];
  _RAND_48 = {1{`RANDOM}};
  __Bi_3_1 = _RAND_48[18:0];
  _RAND_49 = {1{`RANDOM}};
  __Bi_3_2 = _RAND_49[18:0];
  _RAND_50 = {1{`RANDOM}};
  __Bi_3_3 = _RAND_50[18:0];
  _RAND_51 = {1{`RANDOM}};
  __Bi_3_4 = _RAND_51[18:0];
  _RAND_52 = {1{`RANDOM}};
  __Bi_3_5 = _RAND_52[18:0];
  _RAND_53 = {1{`RANDOM}};
  __Bi_5_3 = _RAND_53[18:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Accumu(
  input         clock,
  input         reset,
  input         io_valid_in,
  output        io_valid_out,
  input         io_flag_job,
  input  [36:0] io_in_from_calc8x8_mat_0,
  input  [36:0] io_in_from_calc8x8_mat_1,
  input  [36:0] io_in_from_calc8x8_mat_2,
  input  [36:0] io_in_from_calc8x8_mat_3,
  input  [36:0] io_in_from_calc8x8_mat_4,
  input  [36:0] io_in_from_calc8x8_mat_5,
  input  [36:0] io_in_from_calc8x8_mat_6,
  input  [36:0] io_in_from_calc8x8_mat_7,
  input  [36:0] io_in_from_calc8x8_mat_8,
  input  [36:0] io_in_from_calc8x8_mat_9,
  input  [36:0] io_in_from_calc8x8_mat_10,
  input  [36:0] io_in_from_calc8x8_mat_11,
  input  [36:0] io_in_from_calc8x8_mat_12,
  input  [36:0] io_in_from_calc8x8_mat_13,
  input  [36:0] io_in_from_calc8x8_mat_14,
  input  [36:0] io_in_from_calc8x8_mat_15,
  input  [36:0] io_in_from_calc8x8_mat_16,
  input  [36:0] io_in_from_calc8x8_mat_17,
  input  [36:0] io_in_from_calc8x8_mat_18,
  input  [36:0] io_in_from_calc8x8_mat_19,
  input  [36:0] io_in_from_calc8x8_mat_20,
  input  [36:0] io_in_from_calc8x8_mat_21,
  input  [36:0] io_in_from_calc8x8_mat_22,
  input  [36:0] io_in_from_calc8x8_mat_23,
  input  [36:0] io_in_from_calc8x8_mat_24,
  input  [36:0] io_in_from_calc8x8_mat_25,
  input  [36:0] io_in_from_calc8x8_mat_26,
  input  [36:0] io_in_from_calc8x8_mat_27,
  input  [36:0] io_in_from_calc8x8_mat_28,
  input  [36:0] io_in_from_calc8x8_mat_29,
  input  [36:0] io_in_from_calc8x8_mat_30,
  input  [36:0] io_in_from_calc8x8_mat_31,
  input  [36:0] io_in_from_calc8x8_mat_32,
  input  [36:0] io_in_from_calc8x8_mat_33,
  input  [36:0] io_in_from_calc8x8_mat_34,
  input  [36:0] io_in_from_calc8x8_mat_35,
  input  [36:0] io_in_from_calc8x8_mat_36,
  input  [36:0] io_in_from_calc8x8_mat_37,
  input  [36:0] io_in_from_calc8x8_mat_38,
  input  [36:0] io_in_from_calc8x8_mat_39,
  input  [36:0] io_in_from_calc8x8_mat_40,
  input  [36:0] io_in_from_calc8x8_mat_41,
  input  [36:0] io_in_from_calc8x8_mat_42,
  input  [36:0] io_in_from_calc8x8_mat_43,
  input  [36:0] io_in_from_calc8x8_mat_44,
  input  [36:0] io_in_from_calc8x8_mat_45,
  input  [36:0] io_in_from_calc8x8_mat_46,
  input  [36:0] io_in_from_calc8x8_mat_47,
  input  [36:0] io_in_from_calc8x8_mat_48,
  input  [36:0] io_in_from_calc8x8_mat_49,
  input  [36:0] io_in_from_calc8x8_mat_50,
  input  [36:0] io_in_from_calc8x8_mat_51,
  input  [36:0] io_in_from_calc8x8_mat_52,
  input  [36:0] io_in_from_calc8x8_mat_53,
  input  [36:0] io_in_from_calc8x8_mat_54,
  input  [36:0] io_in_from_calc8x8_mat_55,
  input  [36:0] io_in_from_calc8x8_mat_56,
  input  [36:0] io_in_from_calc8x8_mat_57,
  input  [36:0] io_in_from_calc8x8_mat_58,
  input  [36:0] io_in_from_calc8x8_mat_59,
  input  [36:0] io_in_from_calc8x8_mat_60,
  input  [36:0] io_in_from_calc8x8_mat_61,
  input  [36:0] io_in_from_calc8x8_mat_62,
  input  [36:0] io_in_from_calc8x8_mat_63,
  output [43:0] io_result_mat_0,
  output [43:0] io_result_mat_1,
  output [43:0] io_result_mat_2,
  output [43:0] io_result_mat_3,
  output [43:0] io_result_mat_4,
  output [43:0] io_result_mat_5,
  output [43:0] io_result_mat_6,
  output [43:0] io_result_mat_7,
  output [43:0] io_result_mat_8,
  output [43:0] io_result_mat_9,
  output [43:0] io_result_mat_10,
  output [43:0] io_result_mat_11,
  output [43:0] io_result_mat_12,
  output [43:0] io_result_mat_13,
  output [43:0] io_result_mat_14,
  output [43:0] io_result_mat_15,
  output [43:0] io_result_mat_16,
  output [43:0] io_result_mat_17,
  output [43:0] io_result_mat_18,
  output [43:0] io_result_mat_19,
  output [43:0] io_result_mat_20,
  output [43:0] io_result_mat_21,
  output [43:0] io_result_mat_22,
  output [43:0] io_result_mat_23,
  output [43:0] io_result_mat_24,
  output [43:0] io_result_mat_25,
  output [43:0] io_result_mat_26,
  output [43:0] io_result_mat_27,
  output [43:0] io_result_mat_28,
  output [43:0] io_result_mat_29,
  output [43:0] io_result_mat_30,
  output [43:0] io_result_mat_31,
  output [43:0] io_result_mat_32,
  output [43:0] io_result_mat_33,
  output [43:0] io_result_mat_34,
  output [43:0] io_result_mat_35,
  output [43:0] io_result_mat_36,
  output [43:0] io_result_mat_37,
  output [43:0] io_result_mat_38,
  output [43:0] io_result_mat_39,
  output [43:0] io_result_mat_40,
  output [43:0] io_result_mat_41,
  output [43:0] io_result_mat_42,
  output [43:0] io_result_mat_43,
  output [43:0] io_result_mat_44,
  output [43:0] io_result_mat_45,
  output [43:0] io_result_mat_46,
  output [43:0] io_result_mat_47,
  output [43:0] io_result_mat_48,
  output [43:0] io_result_mat_49,
  output [43:0] io_result_mat_50,
  output [43:0] io_result_mat_51,
  output [43:0] io_result_mat_52,
  output [43:0] io_result_mat_53,
  output [43:0] io_result_mat_54,
  output [43:0] io_result_mat_55,
  output [43:0] io_result_mat_56,
  output [43:0] io_result_mat_57,
  output [43:0] io_result_mat_58,
  output [43:0] io_result_mat_59,
  output [43:0] io_result_mat_60,
  output [43:0] io_result_mat_61,
  output [43:0] io_result_mat_62,
  output [43:0] io_result_mat_63,
  input  [9:0]  io_csum,
  input  [9:0]  io_bias_end_addr,
  output [9:0]  io_bias_addr,
  input  [35:0] io_bias_in,
  input         io_is_in_use
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] counter_ccnt; // @[accumu.scala 27:26]
  reg [9:0] counter_cend; // @[accumu.scala 27:26]
  reg [43:0] output_mat_0; // @[accumu.scala 28:25]
  reg [43:0] output_mat_1; // @[accumu.scala 28:25]
  reg [43:0] output_mat_2; // @[accumu.scala 28:25]
  reg [43:0] output_mat_3; // @[accumu.scala 28:25]
  reg [43:0] output_mat_4; // @[accumu.scala 28:25]
  reg [43:0] output_mat_5; // @[accumu.scala 28:25]
  reg [43:0] output_mat_6; // @[accumu.scala 28:25]
  reg [43:0] output_mat_7; // @[accumu.scala 28:25]
  reg [43:0] output_mat_8; // @[accumu.scala 28:25]
  reg [43:0] output_mat_9; // @[accumu.scala 28:25]
  reg [43:0] output_mat_10; // @[accumu.scala 28:25]
  reg [43:0] output_mat_11; // @[accumu.scala 28:25]
  reg [43:0] output_mat_12; // @[accumu.scala 28:25]
  reg [43:0] output_mat_13; // @[accumu.scala 28:25]
  reg [43:0] output_mat_14; // @[accumu.scala 28:25]
  reg [43:0] output_mat_15; // @[accumu.scala 28:25]
  reg [43:0] output_mat_16; // @[accumu.scala 28:25]
  reg [43:0] output_mat_17; // @[accumu.scala 28:25]
  reg [43:0] output_mat_18; // @[accumu.scala 28:25]
  reg [43:0] output_mat_19; // @[accumu.scala 28:25]
  reg [43:0] output_mat_20; // @[accumu.scala 28:25]
  reg [43:0] output_mat_21; // @[accumu.scala 28:25]
  reg [43:0] output_mat_22; // @[accumu.scala 28:25]
  reg [43:0] output_mat_23; // @[accumu.scala 28:25]
  reg [43:0] output_mat_24; // @[accumu.scala 28:25]
  reg [43:0] output_mat_25; // @[accumu.scala 28:25]
  reg [43:0] output_mat_26; // @[accumu.scala 28:25]
  reg [43:0] output_mat_27; // @[accumu.scala 28:25]
  reg [43:0] output_mat_28; // @[accumu.scala 28:25]
  reg [43:0] output_mat_29; // @[accumu.scala 28:25]
  reg [43:0] output_mat_30; // @[accumu.scala 28:25]
  reg [43:0] output_mat_31; // @[accumu.scala 28:25]
  reg [43:0] output_mat_32; // @[accumu.scala 28:25]
  reg [43:0] output_mat_33; // @[accumu.scala 28:25]
  reg [43:0] output_mat_34; // @[accumu.scala 28:25]
  reg [43:0] output_mat_35; // @[accumu.scala 28:25]
  reg [43:0] output_mat_36; // @[accumu.scala 28:25]
  reg [43:0] output_mat_37; // @[accumu.scala 28:25]
  reg [43:0] output_mat_38; // @[accumu.scala 28:25]
  reg [43:0] output_mat_39; // @[accumu.scala 28:25]
  reg [43:0] output_mat_40; // @[accumu.scala 28:25]
  reg [43:0] output_mat_41; // @[accumu.scala 28:25]
  reg [43:0] output_mat_42; // @[accumu.scala 28:25]
  reg [43:0] output_mat_43; // @[accumu.scala 28:25]
  reg [43:0] output_mat_44; // @[accumu.scala 28:25]
  reg [43:0] output_mat_45; // @[accumu.scala 28:25]
  reg [43:0] output_mat_46; // @[accumu.scala 28:25]
  reg [43:0] output_mat_47; // @[accumu.scala 28:25]
  reg [43:0] output_mat_48; // @[accumu.scala 28:25]
  reg [43:0] output_mat_49; // @[accumu.scala 28:25]
  reg [43:0] output_mat_50; // @[accumu.scala 28:25]
  reg [43:0] output_mat_51; // @[accumu.scala 28:25]
  reg [43:0] output_mat_52; // @[accumu.scala 28:25]
  reg [43:0] output_mat_53; // @[accumu.scala 28:25]
  reg [43:0] output_mat_54; // @[accumu.scala 28:25]
  reg [43:0] output_mat_55; // @[accumu.scala 28:25]
  reg [43:0] output_mat_56; // @[accumu.scala 28:25]
  reg [43:0] output_mat_57; // @[accumu.scala 28:25]
  reg [43:0] output_mat_58; // @[accumu.scala 28:25]
  reg [43:0] output_mat_59; // @[accumu.scala 28:25]
  reg [43:0] output_mat_60; // @[accumu.scala 28:25]
  reg [43:0] output_mat_61; // @[accumu.scala 28:25]
  reg [43:0] output_mat_62; // @[accumu.scala 28:25]
  reg [43:0] output_mat_63; // @[accumu.scala 28:25]
  reg [9:0] now_addr_ccnt; // @[accumu.scala 29:27]
  reg [9:0] now_addr_cend; // @[accumu.scala 29:27]
  reg  enable; // @[accumu.scala 30:25]
  wire [36:0] _GEN_657 = {{1{io_bias_in[35]}},io_bias_in}; // @[accumu.scala 46:63]
  wire [36:0] _output_mat_0_T_2 = $signed(io_in_from_calc8x8_mat_0) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_1_T_2 = $signed(io_in_from_calc8x8_mat_1) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_2_T_2 = $signed(io_in_from_calc8x8_mat_2) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_3_T_2 = $signed(io_in_from_calc8x8_mat_3) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_4_T_2 = $signed(io_in_from_calc8x8_mat_4) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_5_T_2 = $signed(io_in_from_calc8x8_mat_5) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_6_T_2 = $signed(io_in_from_calc8x8_mat_6) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_7_T_2 = $signed(io_in_from_calc8x8_mat_7) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_8_T_2 = $signed(io_in_from_calc8x8_mat_8) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_9_T_2 = $signed(io_in_from_calc8x8_mat_9) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_10_T_2 = $signed(io_in_from_calc8x8_mat_10) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_11_T_2 = $signed(io_in_from_calc8x8_mat_11) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_12_T_2 = $signed(io_in_from_calc8x8_mat_12) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_13_T_2 = $signed(io_in_from_calc8x8_mat_13) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_14_T_2 = $signed(io_in_from_calc8x8_mat_14) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_15_T_2 = $signed(io_in_from_calc8x8_mat_15) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_16_T_2 = $signed(io_in_from_calc8x8_mat_16) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_17_T_2 = $signed(io_in_from_calc8x8_mat_17) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_18_T_2 = $signed(io_in_from_calc8x8_mat_18) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_19_T_2 = $signed(io_in_from_calc8x8_mat_19) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_20_T_2 = $signed(io_in_from_calc8x8_mat_20) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_21_T_2 = $signed(io_in_from_calc8x8_mat_21) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_22_T_2 = $signed(io_in_from_calc8x8_mat_22) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_23_T_2 = $signed(io_in_from_calc8x8_mat_23) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_24_T_2 = $signed(io_in_from_calc8x8_mat_24) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_25_T_2 = $signed(io_in_from_calc8x8_mat_25) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_26_T_2 = $signed(io_in_from_calc8x8_mat_26) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_27_T_2 = $signed(io_in_from_calc8x8_mat_27) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_28_T_2 = $signed(io_in_from_calc8x8_mat_28) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_29_T_2 = $signed(io_in_from_calc8x8_mat_29) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_30_T_2 = $signed(io_in_from_calc8x8_mat_30) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_31_T_2 = $signed(io_in_from_calc8x8_mat_31) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_32_T_2 = $signed(io_in_from_calc8x8_mat_32) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_33_T_2 = $signed(io_in_from_calc8x8_mat_33) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_34_T_2 = $signed(io_in_from_calc8x8_mat_34) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_35_T_2 = $signed(io_in_from_calc8x8_mat_35) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_36_T_2 = $signed(io_in_from_calc8x8_mat_36) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_37_T_2 = $signed(io_in_from_calc8x8_mat_37) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_38_T_2 = $signed(io_in_from_calc8x8_mat_38) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_39_T_2 = $signed(io_in_from_calc8x8_mat_39) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_40_T_2 = $signed(io_in_from_calc8x8_mat_40) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_41_T_2 = $signed(io_in_from_calc8x8_mat_41) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_42_T_2 = $signed(io_in_from_calc8x8_mat_42) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_43_T_2 = $signed(io_in_from_calc8x8_mat_43) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_44_T_2 = $signed(io_in_from_calc8x8_mat_44) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_45_T_2 = $signed(io_in_from_calc8x8_mat_45) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_46_T_2 = $signed(io_in_from_calc8x8_mat_46) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_47_T_2 = $signed(io_in_from_calc8x8_mat_47) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_48_T_2 = $signed(io_in_from_calc8x8_mat_48) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_49_T_2 = $signed(io_in_from_calc8x8_mat_49) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_50_T_2 = $signed(io_in_from_calc8x8_mat_50) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_51_T_2 = $signed(io_in_from_calc8x8_mat_51) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_52_T_2 = $signed(io_in_from_calc8x8_mat_52) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_53_T_2 = $signed(io_in_from_calc8x8_mat_53) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_54_T_2 = $signed(io_in_from_calc8x8_mat_54) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_55_T_2 = $signed(io_in_from_calc8x8_mat_55) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_56_T_2 = $signed(io_in_from_calc8x8_mat_56) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_57_T_2 = $signed(io_in_from_calc8x8_mat_57) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_58_T_2 = $signed(io_in_from_calc8x8_mat_58) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_59_T_2 = $signed(io_in_from_calc8x8_mat_59) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_60_T_2 = $signed(io_in_from_calc8x8_mat_60) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_61_T_2 = $signed(io_in_from_calc8x8_mat_61) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_62_T_2 = $signed(io_in_from_calc8x8_mat_62) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [36:0] _output_mat_63_T_2 = $signed(io_in_from_calc8x8_mat_63) + $signed(_GEN_657); // @[accumu.scala 46:63]
  wire [9:0] _counter_ccnt_T_1 = counter_ccnt - 10'h1; // @[accumu.scala 47:45]
  wire  _T_1 = counter_ccnt == 10'h0; // @[accumu.scala 48:36]
  wire [43:0] _GEN_721 = {{7{io_in_from_calc8x8_mat_0[36]}},io_in_from_calc8x8_mat_0}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_0_T_2 = $signed(_GEN_721) + $signed(output_mat_0); // @[accumu.scala 51:66]
  wire [43:0] _GEN_722 = {{7{io_in_from_calc8x8_mat_1[36]}},io_in_from_calc8x8_mat_1}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_1_T_2 = $signed(_GEN_722) + $signed(output_mat_1); // @[accumu.scala 51:66]
  wire [43:0] _GEN_723 = {{7{io_in_from_calc8x8_mat_2[36]}},io_in_from_calc8x8_mat_2}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_2_T_2 = $signed(_GEN_723) + $signed(output_mat_2); // @[accumu.scala 51:66]
  wire [43:0] _GEN_724 = {{7{io_in_from_calc8x8_mat_3[36]}},io_in_from_calc8x8_mat_3}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_3_T_2 = $signed(_GEN_724) + $signed(output_mat_3); // @[accumu.scala 51:66]
  wire [43:0] _GEN_725 = {{7{io_in_from_calc8x8_mat_4[36]}},io_in_from_calc8x8_mat_4}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_4_T_2 = $signed(_GEN_725) + $signed(output_mat_4); // @[accumu.scala 51:66]
  wire [43:0] _GEN_726 = {{7{io_in_from_calc8x8_mat_5[36]}},io_in_from_calc8x8_mat_5}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_5_T_2 = $signed(_GEN_726) + $signed(output_mat_5); // @[accumu.scala 51:66]
  wire [43:0] _GEN_727 = {{7{io_in_from_calc8x8_mat_6[36]}},io_in_from_calc8x8_mat_6}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_6_T_2 = $signed(_GEN_727) + $signed(output_mat_6); // @[accumu.scala 51:66]
  wire [43:0] _GEN_728 = {{7{io_in_from_calc8x8_mat_7[36]}},io_in_from_calc8x8_mat_7}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_7_T_2 = $signed(_GEN_728) + $signed(output_mat_7); // @[accumu.scala 51:66]
  wire [43:0] _GEN_729 = {{7{io_in_from_calc8x8_mat_8[36]}},io_in_from_calc8x8_mat_8}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_8_T_2 = $signed(_GEN_729) + $signed(output_mat_8); // @[accumu.scala 51:66]
  wire [43:0] _GEN_730 = {{7{io_in_from_calc8x8_mat_9[36]}},io_in_from_calc8x8_mat_9}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_9_T_2 = $signed(_GEN_730) + $signed(output_mat_9); // @[accumu.scala 51:66]
  wire [43:0] _GEN_731 = {{7{io_in_from_calc8x8_mat_10[36]}},io_in_from_calc8x8_mat_10}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_10_T_2 = $signed(_GEN_731) + $signed(output_mat_10); // @[accumu.scala 51:66]
  wire [43:0] _GEN_732 = {{7{io_in_from_calc8x8_mat_11[36]}},io_in_from_calc8x8_mat_11}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_11_T_2 = $signed(_GEN_732) + $signed(output_mat_11); // @[accumu.scala 51:66]
  wire [43:0] _GEN_733 = {{7{io_in_from_calc8x8_mat_12[36]}},io_in_from_calc8x8_mat_12}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_12_T_2 = $signed(_GEN_733) + $signed(output_mat_12); // @[accumu.scala 51:66]
  wire [43:0] _GEN_734 = {{7{io_in_from_calc8x8_mat_13[36]}},io_in_from_calc8x8_mat_13}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_13_T_2 = $signed(_GEN_734) + $signed(output_mat_13); // @[accumu.scala 51:66]
  wire [43:0] _GEN_735 = {{7{io_in_from_calc8x8_mat_14[36]}},io_in_from_calc8x8_mat_14}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_14_T_2 = $signed(_GEN_735) + $signed(output_mat_14); // @[accumu.scala 51:66]
  wire [43:0] _GEN_736 = {{7{io_in_from_calc8x8_mat_15[36]}},io_in_from_calc8x8_mat_15}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_15_T_2 = $signed(_GEN_736) + $signed(output_mat_15); // @[accumu.scala 51:66]
  wire [43:0] _GEN_737 = {{7{io_in_from_calc8x8_mat_16[36]}},io_in_from_calc8x8_mat_16}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_16_T_2 = $signed(_GEN_737) + $signed(output_mat_16); // @[accumu.scala 51:66]
  wire [43:0] _GEN_738 = {{7{io_in_from_calc8x8_mat_17[36]}},io_in_from_calc8x8_mat_17}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_17_T_2 = $signed(_GEN_738) + $signed(output_mat_17); // @[accumu.scala 51:66]
  wire [43:0] _GEN_739 = {{7{io_in_from_calc8x8_mat_18[36]}},io_in_from_calc8x8_mat_18}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_18_T_2 = $signed(_GEN_739) + $signed(output_mat_18); // @[accumu.scala 51:66]
  wire [43:0] _GEN_740 = {{7{io_in_from_calc8x8_mat_19[36]}},io_in_from_calc8x8_mat_19}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_19_T_2 = $signed(_GEN_740) + $signed(output_mat_19); // @[accumu.scala 51:66]
  wire [43:0] _GEN_741 = {{7{io_in_from_calc8x8_mat_20[36]}},io_in_from_calc8x8_mat_20}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_20_T_2 = $signed(_GEN_741) + $signed(output_mat_20); // @[accumu.scala 51:66]
  wire [43:0] _GEN_742 = {{7{io_in_from_calc8x8_mat_21[36]}},io_in_from_calc8x8_mat_21}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_21_T_2 = $signed(_GEN_742) + $signed(output_mat_21); // @[accumu.scala 51:66]
  wire [43:0] _GEN_743 = {{7{io_in_from_calc8x8_mat_22[36]}},io_in_from_calc8x8_mat_22}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_22_T_2 = $signed(_GEN_743) + $signed(output_mat_22); // @[accumu.scala 51:66]
  wire [43:0] _GEN_744 = {{7{io_in_from_calc8x8_mat_23[36]}},io_in_from_calc8x8_mat_23}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_23_T_2 = $signed(_GEN_744) + $signed(output_mat_23); // @[accumu.scala 51:66]
  wire [43:0] _GEN_745 = {{7{io_in_from_calc8x8_mat_24[36]}},io_in_from_calc8x8_mat_24}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_24_T_2 = $signed(_GEN_745) + $signed(output_mat_24); // @[accumu.scala 51:66]
  wire [43:0] _GEN_746 = {{7{io_in_from_calc8x8_mat_25[36]}},io_in_from_calc8x8_mat_25}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_25_T_2 = $signed(_GEN_746) + $signed(output_mat_25); // @[accumu.scala 51:66]
  wire [43:0] _GEN_747 = {{7{io_in_from_calc8x8_mat_26[36]}},io_in_from_calc8x8_mat_26}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_26_T_2 = $signed(_GEN_747) + $signed(output_mat_26); // @[accumu.scala 51:66]
  wire [43:0] _GEN_748 = {{7{io_in_from_calc8x8_mat_27[36]}},io_in_from_calc8x8_mat_27}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_27_T_2 = $signed(_GEN_748) + $signed(output_mat_27); // @[accumu.scala 51:66]
  wire [43:0] _GEN_749 = {{7{io_in_from_calc8x8_mat_28[36]}},io_in_from_calc8x8_mat_28}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_28_T_2 = $signed(_GEN_749) + $signed(output_mat_28); // @[accumu.scala 51:66]
  wire [43:0] _GEN_750 = {{7{io_in_from_calc8x8_mat_29[36]}},io_in_from_calc8x8_mat_29}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_29_T_2 = $signed(_GEN_750) + $signed(output_mat_29); // @[accumu.scala 51:66]
  wire [43:0] _GEN_751 = {{7{io_in_from_calc8x8_mat_30[36]}},io_in_from_calc8x8_mat_30}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_30_T_2 = $signed(_GEN_751) + $signed(output_mat_30); // @[accumu.scala 51:66]
  wire [43:0] _GEN_752 = {{7{io_in_from_calc8x8_mat_31[36]}},io_in_from_calc8x8_mat_31}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_31_T_2 = $signed(_GEN_752) + $signed(output_mat_31); // @[accumu.scala 51:66]
  wire [43:0] _GEN_753 = {{7{io_in_from_calc8x8_mat_32[36]}},io_in_from_calc8x8_mat_32}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_32_T_2 = $signed(_GEN_753) + $signed(output_mat_32); // @[accumu.scala 51:66]
  wire [43:0] _GEN_754 = {{7{io_in_from_calc8x8_mat_33[36]}},io_in_from_calc8x8_mat_33}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_33_T_2 = $signed(_GEN_754) + $signed(output_mat_33); // @[accumu.scala 51:66]
  wire [43:0] _GEN_755 = {{7{io_in_from_calc8x8_mat_34[36]}},io_in_from_calc8x8_mat_34}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_34_T_2 = $signed(_GEN_755) + $signed(output_mat_34); // @[accumu.scala 51:66]
  wire [43:0] _GEN_756 = {{7{io_in_from_calc8x8_mat_35[36]}},io_in_from_calc8x8_mat_35}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_35_T_2 = $signed(_GEN_756) + $signed(output_mat_35); // @[accumu.scala 51:66]
  wire [43:0] _GEN_757 = {{7{io_in_from_calc8x8_mat_36[36]}},io_in_from_calc8x8_mat_36}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_36_T_2 = $signed(_GEN_757) + $signed(output_mat_36); // @[accumu.scala 51:66]
  wire [43:0] _GEN_758 = {{7{io_in_from_calc8x8_mat_37[36]}},io_in_from_calc8x8_mat_37}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_37_T_2 = $signed(_GEN_758) + $signed(output_mat_37); // @[accumu.scala 51:66]
  wire [43:0] _GEN_759 = {{7{io_in_from_calc8x8_mat_38[36]}},io_in_from_calc8x8_mat_38}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_38_T_2 = $signed(_GEN_759) + $signed(output_mat_38); // @[accumu.scala 51:66]
  wire [43:0] _GEN_760 = {{7{io_in_from_calc8x8_mat_39[36]}},io_in_from_calc8x8_mat_39}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_39_T_2 = $signed(_GEN_760) + $signed(output_mat_39); // @[accumu.scala 51:66]
  wire [43:0] _GEN_761 = {{7{io_in_from_calc8x8_mat_40[36]}},io_in_from_calc8x8_mat_40}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_40_T_2 = $signed(_GEN_761) + $signed(output_mat_40); // @[accumu.scala 51:66]
  wire [43:0] _GEN_762 = {{7{io_in_from_calc8x8_mat_41[36]}},io_in_from_calc8x8_mat_41}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_41_T_2 = $signed(_GEN_762) + $signed(output_mat_41); // @[accumu.scala 51:66]
  wire [43:0] _GEN_763 = {{7{io_in_from_calc8x8_mat_42[36]}},io_in_from_calc8x8_mat_42}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_42_T_2 = $signed(_GEN_763) + $signed(output_mat_42); // @[accumu.scala 51:66]
  wire [43:0] _GEN_764 = {{7{io_in_from_calc8x8_mat_43[36]}},io_in_from_calc8x8_mat_43}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_43_T_2 = $signed(_GEN_764) + $signed(output_mat_43); // @[accumu.scala 51:66]
  wire [43:0] _GEN_765 = {{7{io_in_from_calc8x8_mat_44[36]}},io_in_from_calc8x8_mat_44}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_44_T_2 = $signed(_GEN_765) + $signed(output_mat_44); // @[accumu.scala 51:66]
  wire [43:0] _GEN_766 = {{7{io_in_from_calc8x8_mat_45[36]}},io_in_from_calc8x8_mat_45}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_45_T_2 = $signed(_GEN_766) + $signed(output_mat_45); // @[accumu.scala 51:66]
  wire [43:0] _GEN_767 = {{7{io_in_from_calc8x8_mat_46[36]}},io_in_from_calc8x8_mat_46}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_46_T_2 = $signed(_GEN_767) + $signed(output_mat_46); // @[accumu.scala 51:66]
  wire [43:0] _GEN_768 = {{7{io_in_from_calc8x8_mat_47[36]}},io_in_from_calc8x8_mat_47}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_47_T_2 = $signed(_GEN_768) + $signed(output_mat_47); // @[accumu.scala 51:66]
  wire [43:0] _GEN_769 = {{7{io_in_from_calc8x8_mat_48[36]}},io_in_from_calc8x8_mat_48}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_48_T_2 = $signed(_GEN_769) + $signed(output_mat_48); // @[accumu.scala 51:66]
  wire [43:0] _GEN_770 = {{7{io_in_from_calc8x8_mat_49[36]}},io_in_from_calc8x8_mat_49}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_49_T_2 = $signed(_GEN_770) + $signed(output_mat_49); // @[accumu.scala 51:66]
  wire [43:0] _GEN_771 = {{7{io_in_from_calc8x8_mat_50[36]}},io_in_from_calc8x8_mat_50}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_50_T_2 = $signed(_GEN_771) + $signed(output_mat_50); // @[accumu.scala 51:66]
  wire [43:0] _GEN_772 = {{7{io_in_from_calc8x8_mat_51[36]}},io_in_from_calc8x8_mat_51}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_51_T_2 = $signed(_GEN_772) + $signed(output_mat_51); // @[accumu.scala 51:66]
  wire [43:0] _GEN_773 = {{7{io_in_from_calc8x8_mat_52[36]}},io_in_from_calc8x8_mat_52}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_52_T_2 = $signed(_GEN_773) + $signed(output_mat_52); // @[accumu.scala 51:66]
  wire [43:0] _GEN_774 = {{7{io_in_from_calc8x8_mat_53[36]}},io_in_from_calc8x8_mat_53}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_53_T_2 = $signed(_GEN_774) + $signed(output_mat_53); // @[accumu.scala 51:66]
  wire [43:0] _GEN_775 = {{7{io_in_from_calc8x8_mat_54[36]}},io_in_from_calc8x8_mat_54}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_54_T_2 = $signed(_GEN_775) + $signed(output_mat_54); // @[accumu.scala 51:66]
  wire [43:0] _GEN_776 = {{7{io_in_from_calc8x8_mat_55[36]}},io_in_from_calc8x8_mat_55}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_55_T_2 = $signed(_GEN_776) + $signed(output_mat_55); // @[accumu.scala 51:66]
  wire [43:0] _GEN_777 = {{7{io_in_from_calc8x8_mat_56[36]}},io_in_from_calc8x8_mat_56}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_56_T_2 = $signed(_GEN_777) + $signed(output_mat_56); // @[accumu.scala 51:66]
  wire [43:0] _GEN_778 = {{7{io_in_from_calc8x8_mat_57[36]}},io_in_from_calc8x8_mat_57}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_57_T_2 = $signed(_GEN_778) + $signed(output_mat_57); // @[accumu.scala 51:66]
  wire [43:0] _GEN_779 = {{7{io_in_from_calc8x8_mat_58[36]}},io_in_from_calc8x8_mat_58}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_58_T_2 = $signed(_GEN_779) + $signed(output_mat_58); // @[accumu.scala 51:66]
  wire [43:0] _GEN_780 = {{7{io_in_from_calc8x8_mat_59[36]}},io_in_from_calc8x8_mat_59}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_59_T_2 = $signed(_GEN_780) + $signed(output_mat_59); // @[accumu.scala 51:66]
  wire [43:0] _GEN_781 = {{7{io_in_from_calc8x8_mat_60[36]}},io_in_from_calc8x8_mat_60}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_60_T_2 = $signed(_GEN_781) + $signed(output_mat_60); // @[accumu.scala 51:66]
  wire [43:0] _GEN_782 = {{7{io_in_from_calc8x8_mat_61[36]}},io_in_from_calc8x8_mat_61}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_61_T_2 = $signed(_GEN_782) + $signed(output_mat_61); // @[accumu.scala 51:66]
  wire [43:0] _GEN_783 = {{7{io_in_from_calc8x8_mat_62[36]}},io_in_from_calc8x8_mat_62}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_62_T_2 = $signed(_GEN_783) + $signed(output_mat_62); // @[accumu.scala 51:66]
  wire [43:0] _GEN_784 = {{7{io_in_from_calc8x8_mat_63[36]}},io_in_from_calc8x8_mat_63}; // @[accumu.scala 51:66]
  wire [43:0] _io_result_mat_63_T_2 = $signed(_GEN_784) + $signed(output_mat_63); // @[accumu.scala 51:66]
  wire [43:0] _output_mat_0_T_5 = $signed(output_mat_0) + $signed(_GEN_721); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_1_T_5 = $signed(output_mat_1) + $signed(_GEN_722); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_2_T_5 = $signed(output_mat_2) + $signed(_GEN_723); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_3_T_5 = $signed(output_mat_3) + $signed(_GEN_724); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_4_T_5 = $signed(output_mat_4) + $signed(_GEN_725); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_5_T_5 = $signed(output_mat_5) + $signed(_GEN_726); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_6_T_5 = $signed(output_mat_6) + $signed(_GEN_727); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_7_T_5 = $signed(output_mat_7) + $signed(_GEN_728); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_8_T_5 = $signed(output_mat_8) + $signed(_GEN_729); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_9_T_5 = $signed(output_mat_9) + $signed(_GEN_730); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_10_T_5 = $signed(output_mat_10) + $signed(_GEN_731); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_11_T_5 = $signed(output_mat_11) + $signed(_GEN_732); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_12_T_5 = $signed(output_mat_12) + $signed(_GEN_733); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_13_T_5 = $signed(output_mat_13) + $signed(_GEN_734); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_14_T_5 = $signed(output_mat_14) + $signed(_GEN_735); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_15_T_5 = $signed(output_mat_15) + $signed(_GEN_736); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_16_T_5 = $signed(output_mat_16) + $signed(_GEN_737); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_17_T_5 = $signed(output_mat_17) + $signed(_GEN_738); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_18_T_5 = $signed(output_mat_18) + $signed(_GEN_739); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_19_T_5 = $signed(output_mat_19) + $signed(_GEN_740); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_20_T_5 = $signed(output_mat_20) + $signed(_GEN_741); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_21_T_5 = $signed(output_mat_21) + $signed(_GEN_742); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_22_T_5 = $signed(output_mat_22) + $signed(_GEN_743); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_23_T_5 = $signed(output_mat_23) + $signed(_GEN_744); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_24_T_5 = $signed(output_mat_24) + $signed(_GEN_745); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_25_T_5 = $signed(output_mat_25) + $signed(_GEN_746); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_26_T_5 = $signed(output_mat_26) + $signed(_GEN_747); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_27_T_5 = $signed(output_mat_27) + $signed(_GEN_748); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_28_T_5 = $signed(output_mat_28) + $signed(_GEN_749); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_29_T_5 = $signed(output_mat_29) + $signed(_GEN_750); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_30_T_5 = $signed(output_mat_30) + $signed(_GEN_751); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_31_T_5 = $signed(output_mat_31) + $signed(_GEN_752); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_32_T_5 = $signed(output_mat_32) + $signed(_GEN_753); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_33_T_5 = $signed(output_mat_33) + $signed(_GEN_754); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_34_T_5 = $signed(output_mat_34) + $signed(_GEN_755); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_35_T_5 = $signed(output_mat_35) + $signed(_GEN_756); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_36_T_5 = $signed(output_mat_36) + $signed(_GEN_757); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_37_T_5 = $signed(output_mat_37) + $signed(_GEN_758); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_38_T_5 = $signed(output_mat_38) + $signed(_GEN_759); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_39_T_5 = $signed(output_mat_39) + $signed(_GEN_760); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_40_T_5 = $signed(output_mat_40) + $signed(_GEN_761); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_41_T_5 = $signed(output_mat_41) + $signed(_GEN_762); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_42_T_5 = $signed(output_mat_42) + $signed(_GEN_763); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_43_T_5 = $signed(output_mat_43) + $signed(_GEN_764); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_44_T_5 = $signed(output_mat_44) + $signed(_GEN_765); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_45_T_5 = $signed(output_mat_45) + $signed(_GEN_766); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_46_T_5 = $signed(output_mat_46) + $signed(_GEN_767); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_47_T_5 = $signed(output_mat_47) + $signed(_GEN_768); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_48_T_5 = $signed(output_mat_48) + $signed(_GEN_769); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_49_T_5 = $signed(output_mat_49) + $signed(_GEN_770); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_50_T_5 = $signed(output_mat_50) + $signed(_GEN_771); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_51_T_5 = $signed(output_mat_51) + $signed(_GEN_772); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_52_T_5 = $signed(output_mat_52) + $signed(_GEN_773); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_53_T_5 = $signed(output_mat_53) + $signed(_GEN_774); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_54_T_5 = $signed(output_mat_54) + $signed(_GEN_775); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_55_T_5 = $signed(output_mat_55) + $signed(_GEN_776); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_56_T_5 = $signed(output_mat_56) + $signed(_GEN_777); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_57_T_5 = $signed(output_mat_57) + $signed(_GEN_778); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_58_T_5 = $signed(output_mat_58) + $signed(_GEN_779); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_59_T_5 = $signed(output_mat_59) + $signed(_GEN_780); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_60_T_5 = $signed(output_mat_60) + $signed(_GEN_781); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_61_T_5 = $signed(output_mat_61) + $signed(_GEN_782); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_62_T_5 = $signed(output_mat_62) + $signed(_GEN_783); // @[accumu.scala 56:51]
  wire [43:0] _output_mat_63_T_5 = $signed(output_mat_63) + $signed(_GEN_784); // @[accumu.scala 56:51]
  wire [43:0] _GEN_1 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_0_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_2 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_1_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_3 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_2_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_4 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_3_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_5 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_4_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_6 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_5_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_7 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_6_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_8 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_7_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_9 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_8_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_10 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_9_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_11 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_10_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_12 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_11_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_13 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_12_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_14 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_13_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_15 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_14_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_16 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_15_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_17 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_16_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_18 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_17_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_19 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_18_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_20 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_19_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_21 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_20_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_22 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_21_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_23 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_22_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_24 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_23_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_25 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_24_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_26 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_25_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_27 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_26_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_28 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_27_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_29 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_28_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_30 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_29_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_31 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_30_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_32 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_31_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_33 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_32_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_34 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_33_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_35 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_34_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_36 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_35_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_37 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_36_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_38 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_37_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_39 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_38_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_40 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_39_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_41 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_40_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_42 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_41_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_43 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_42_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_44 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_43_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_45 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_44_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_46 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_45_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_47 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_46_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_48 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_47_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_49 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_48_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_50 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_49_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_51 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_50_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_52 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_51_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_53 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_52_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_54 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_53_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_55 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_54_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_56 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_55_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_57 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_56_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_58 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_57_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_59 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_58_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_60 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_59_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_61 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_60_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_62 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_61_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_63 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_62_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [43:0] _GEN_64 = counter_ccnt == 10'h0 ? $signed(_io_result_mat_63_T_2) : $signed(44'sh0); // @[accumu.scala 48:43 accumu.scala 51:38 accumu.scala 32:15]
  wire [9:0] _GEN_65 = counter_ccnt == 10'h0 ? counter_cend : _counter_ccnt_T_1; // @[accumu.scala 48:43 accumu.scala 52:30 accumu.scala 57:30]
  wire [43:0] _GEN_66 = counter_ccnt == 10'h0 ? $signed(output_mat_0) : $signed(_output_mat_0_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_67 = counter_ccnt == 10'h0 ? $signed(output_mat_1) : $signed(_output_mat_1_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_68 = counter_ccnt == 10'h0 ? $signed(output_mat_2) : $signed(_output_mat_2_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_69 = counter_ccnt == 10'h0 ? $signed(output_mat_3) : $signed(_output_mat_3_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_70 = counter_ccnt == 10'h0 ? $signed(output_mat_4) : $signed(_output_mat_4_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_71 = counter_ccnt == 10'h0 ? $signed(output_mat_5) : $signed(_output_mat_5_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_72 = counter_ccnt == 10'h0 ? $signed(output_mat_6) : $signed(_output_mat_6_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_73 = counter_ccnt == 10'h0 ? $signed(output_mat_7) : $signed(_output_mat_7_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_74 = counter_ccnt == 10'h0 ? $signed(output_mat_8) : $signed(_output_mat_8_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_75 = counter_ccnt == 10'h0 ? $signed(output_mat_9) : $signed(_output_mat_9_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_76 = counter_ccnt == 10'h0 ? $signed(output_mat_10) : $signed(_output_mat_10_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_77 = counter_ccnt == 10'h0 ? $signed(output_mat_11) : $signed(_output_mat_11_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_78 = counter_ccnt == 10'h0 ? $signed(output_mat_12) : $signed(_output_mat_12_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_79 = counter_ccnt == 10'h0 ? $signed(output_mat_13) : $signed(_output_mat_13_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_80 = counter_ccnt == 10'h0 ? $signed(output_mat_14) : $signed(_output_mat_14_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_81 = counter_ccnt == 10'h0 ? $signed(output_mat_15) : $signed(_output_mat_15_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_82 = counter_ccnt == 10'h0 ? $signed(output_mat_16) : $signed(_output_mat_16_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_83 = counter_ccnt == 10'h0 ? $signed(output_mat_17) : $signed(_output_mat_17_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_84 = counter_ccnt == 10'h0 ? $signed(output_mat_18) : $signed(_output_mat_18_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_85 = counter_ccnt == 10'h0 ? $signed(output_mat_19) : $signed(_output_mat_19_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_86 = counter_ccnt == 10'h0 ? $signed(output_mat_20) : $signed(_output_mat_20_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_87 = counter_ccnt == 10'h0 ? $signed(output_mat_21) : $signed(_output_mat_21_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_88 = counter_ccnt == 10'h0 ? $signed(output_mat_22) : $signed(_output_mat_22_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_89 = counter_ccnt == 10'h0 ? $signed(output_mat_23) : $signed(_output_mat_23_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_90 = counter_ccnt == 10'h0 ? $signed(output_mat_24) : $signed(_output_mat_24_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_91 = counter_ccnt == 10'h0 ? $signed(output_mat_25) : $signed(_output_mat_25_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_92 = counter_ccnt == 10'h0 ? $signed(output_mat_26) : $signed(_output_mat_26_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_93 = counter_ccnt == 10'h0 ? $signed(output_mat_27) : $signed(_output_mat_27_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_94 = counter_ccnt == 10'h0 ? $signed(output_mat_28) : $signed(_output_mat_28_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_95 = counter_ccnt == 10'h0 ? $signed(output_mat_29) : $signed(_output_mat_29_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_96 = counter_ccnt == 10'h0 ? $signed(output_mat_30) : $signed(_output_mat_30_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_97 = counter_ccnt == 10'h0 ? $signed(output_mat_31) : $signed(_output_mat_31_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_98 = counter_ccnt == 10'h0 ? $signed(output_mat_32) : $signed(_output_mat_32_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_99 = counter_ccnt == 10'h0 ? $signed(output_mat_33) : $signed(_output_mat_33_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_100 = counter_ccnt == 10'h0 ? $signed(output_mat_34) : $signed(_output_mat_34_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_101 = counter_ccnt == 10'h0 ? $signed(output_mat_35) : $signed(_output_mat_35_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_102 = counter_ccnt == 10'h0 ? $signed(output_mat_36) : $signed(_output_mat_36_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_103 = counter_ccnt == 10'h0 ? $signed(output_mat_37) : $signed(_output_mat_37_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_104 = counter_ccnt == 10'h0 ? $signed(output_mat_38) : $signed(_output_mat_38_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_105 = counter_ccnt == 10'h0 ? $signed(output_mat_39) : $signed(_output_mat_39_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_106 = counter_ccnt == 10'h0 ? $signed(output_mat_40) : $signed(_output_mat_40_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_107 = counter_ccnt == 10'h0 ? $signed(output_mat_41) : $signed(_output_mat_41_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_108 = counter_ccnt == 10'h0 ? $signed(output_mat_42) : $signed(_output_mat_42_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_109 = counter_ccnt == 10'h0 ? $signed(output_mat_43) : $signed(_output_mat_43_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_110 = counter_ccnt == 10'h0 ? $signed(output_mat_44) : $signed(_output_mat_44_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_111 = counter_ccnt == 10'h0 ? $signed(output_mat_45) : $signed(_output_mat_45_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_112 = counter_ccnt == 10'h0 ? $signed(output_mat_46) : $signed(_output_mat_46_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_113 = counter_ccnt == 10'h0 ? $signed(output_mat_47) : $signed(_output_mat_47_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_114 = counter_ccnt == 10'h0 ? $signed(output_mat_48) : $signed(_output_mat_48_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_115 = counter_ccnt == 10'h0 ? $signed(output_mat_49) : $signed(_output_mat_49_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_116 = counter_ccnt == 10'h0 ? $signed(output_mat_50) : $signed(_output_mat_50_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_117 = counter_ccnt == 10'h0 ? $signed(output_mat_51) : $signed(_output_mat_51_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_118 = counter_ccnt == 10'h0 ? $signed(output_mat_52) : $signed(_output_mat_52_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_119 = counter_ccnt == 10'h0 ? $signed(output_mat_53) : $signed(_output_mat_53_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_120 = counter_ccnt == 10'h0 ? $signed(output_mat_54) : $signed(_output_mat_54_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_121 = counter_ccnt == 10'h0 ? $signed(output_mat_55) : $signed(_output_mat_55_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_122 = counter_ccnt == 10'h0 ? $signed(output_mat_56) : $signed(_output_mat_56_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_123 = counter_ccnt == 10'h0 ? $signed(output_mat_57) : $signed(_output_mat_57_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_124 = counter_ccnt == 10'h0 ? $signed(output_mat_58) : $signed(_output_mat_58_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_125 = counter_ccnt == 10'h0 ? $signed(output_mat_59) : $signed(_output_mat_59_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_126 = counter_ccnt == 10'h0 ? $signed(output_mat_60) : $signed(_output_mat_60_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_127 = counter_ccnt == 10'h0 ? $signed(output_mat_61) : $signed(_output_mat_61_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_128 = counter_ccnt == 10'h0 ? $signed(output_mat_62) : $signed(_output_mat_62_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire [43:0] _GEN_129 = counter_ccnt == 10'h0 ? $signed(output_mat_63) : $signed(_output_mat_63_T_5); // @[accumu.scala 48:43 accumu.scala 28:25 accumu.scala 56:35]
  wire  _GEN_130 = counter_ccnt == counter_cend ? 1'h0 : _T_1; // @[accumu.scala 43:46 accumu.scala 44:30]
  wire [43:0] _GEN_131 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_0_T_2[36]}},_output_mat_0_T_2}) :
    $signed(_GEN_66); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_132 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_1_T_2[36]}},_output_mat_1_T_2}) :
    $signed(_GEN_67); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_133 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_2_T_2[36]}},_output_mat_2_T_2}) :
    $signed(_GEN_68); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_134 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_3_T_2[36]}},_output_mat_3_T_2}) :
    $signed(_GEN_69); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_135 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_4_T_2[36]}},_output_mat_4_T_2}) :
    $signed(_GEN_70); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_136 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_5_T_2[36]}},_output_mat_5_T_2}) :
    $signed(_GEN_71); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_137 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_6_T_2[36]}},_output_mat_6_T_2}) :
    $signed(_GEN_72); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_138 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_7_T_2[36]}},_output_mat_7_T_2}) :
    $signed(_GEN_73); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_139 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_8_T_2[36]}},_output_mat_8_T_2}) :
    $signed(_GEN_74); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_140 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_9_T_2[36]}},_output_mat_9_T_2}) :
    $signed(_GEN_75); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_141 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_10_T_2[36]}},_output_mat_10_T_2}) :
    $signed(_GEN_76); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_142 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_11_T_2[36]}},_output_mat_11_T_2}) :
    $signed(_GEN_77); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_143 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_12_T_2[36]}},_output_mat_12_T_2}) :
    $signed(_GEN_78); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_144 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_13_T_2[36]}},_output_mat_13_T_2}) :
    $signed(_GEN_79); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_145 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_14_T_2[36]}},_output_mat_14_T_2}) :
    $signed(_GEN_80); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_146 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_15_T_2[36]}},_output_mat_15_T_2}) :
    $signed(_GEN_81); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_147 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_16_T_2[36]}},_output_mat_16_T_2}) :
    $signed(_GEN_82); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_148 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_17_T_2[36]}},_output_mat_17_T_2}) :
    $signed(_GEN_83); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_149 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_18_T_2[36]}},_output_mat_18_T_2}) :
    $signed(_GEN_84); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_150 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_19_T_2[36]}},_output_mat_19_T_2}) :
    $signed(_GEN_85); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_151 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_20_T_2[36]}},_output_mat_20_T_2}) :
    $signed(_GEN_86); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_152 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_21_T_2[36]}},_output_mat_21_T_2}) :
    $signed(_GEN_87); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_153 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_22_T_2[36]}},_output_mat_22_T_2}) :
    $signed(_GEN_88); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_154 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_23_T_2[36]}},_output_mat_23_T_2}) :
    $signed(_GEN_89); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_155 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_24_T_2[36]}},_output_mat_24_T_2}) :
    $signed(_GEN_90); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_156 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_25_T_2[36]}},_output_mat_25_T_2}) :
    $signed(_GEN_91); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_157 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_26_T_2[36]}},_output_mat_26_T_2}) :
    $signed(_GEN_92); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_158 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_27_T_2[36]}},_output_mat_27_T_2}) :
    $signed(_GEN_93); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_159 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_28_T_2[36]}},_output_mat_28_T_2}) :
    $signed(_GEN_94); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_160 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_29_T_2[36]}},_output_mat_29_T_2}) :
    $signed(_GEN_95); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_161 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_30_T_2[36]}},_output_mat_30_T_2}) :
    $signed(_GEN_96); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_162 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_31_T_2[36]}},_output_mat_31_T_2}) :
    $signed(_GEN_97); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_163 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_32_T_2[36]}},_output_mat_32_T_2}) :
    $signed(_GEN_98); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_164 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_33_T_2[36]}},_output_mat_33_T_2}) :
    $signed(_GEN_99); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_165 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_34_T_2[36]}},_output_mat_34_T_2}) :
    $signed(_GEN_100); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_166 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_35_T_2[36]}},_output_mat_35_T_2}) :
    $signed(_GEN_101); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_167 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_36_T_2[36]}},_output_mat_36_T_2}) :
    $signed(_GEN_102); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_168 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_37_T_2[36]}},_output_mat_37_T_2}) :
    $signed(_GEN_103); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_169 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_38_T_2[36]}},_output_mat_38_T_2}) :
    $signed(_GEN_104); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_170 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_39_T_2[36]}},_output_mat_39_T_2}) :
    $signed(_GEN_105); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_171 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_40_T_2[36]}},_output_mat_40_T_2}) :
    $signed(_GEN_106); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_172 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_41_T_2[36]}},_output_mat_41_T_2}) :
    $signed(_GEN_107); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_173 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_42_T_2[36]}},_output_mat_42_T_2}) :
    $signed(_GEN_108); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_174 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_43_T_2[36]}},_output_mat_43_T_2}) :
    $signed(_GEN_109); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_175 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_44_T_2[36]}},_output_mat_44_T_2}) :
    $signed(_GEN_110); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_176 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_45_T_2[36]}},_output_mat_45_T_2}) :
    $signed(_GEN_111); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_177 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_46_T_2[36]}},_output_mat_46_T_2}) :
    $signed(_GEN_112); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_178 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_47_T_2[36]}},_output_mat_47_T_2}) :
    $signed(_GEN_113); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_179 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_48_T_2[36]}},_output_mat_48_T_2}) :
    $signed(_GEN_114); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_180 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_49_T_2[36]}},_output_mat_49_T_2}) :
    $signed(_GEN_115); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_181 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_50_T_2[36]}},_output_mat_50_T_2}) :
    $signed(_GEN_116); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_182 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_51_T_2[36]}},_output_mat_51_T_2}) :
    $signed(_GEN_117); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_183 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_52_T_2[36]}},_output_mat_52_T_2}) :
    $signed(_GEN_118); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_184 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_53_T_2[36]}},_output_mat_53_T_2}) :
    $signed(_GEN_119); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_185 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_54_T_2[36]}},_output_mat_54_T_2}) :
    $signed(_GEN_120); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_186 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_55_T_2[36]}},_output_mat_55_T_2}) :
    $signed(_GEN_121); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_187 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_56_T_2[36]}},_output_mat_56_T_2}) :
    $signed(_GEN_122); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_188 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_57_T_2[36]}},_output_mat_57_T_2}) :
    $signed(_GEN_123); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_189 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_58_T_2[36]}},_output_mat_58_T_2}) :
    $signed(_GEN_124); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_190 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_59_T_2[36]}},_output_mat_59_T_2}) :
    $signed(_GEN_125); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_191 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_60_T_2[36]}},_output_mat_60_T_2}) :
    $signed(_GEN_126); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_192 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_61_T_2[36]}},_output_mat_61_T_2}) :
    $signed(_GEN_127); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_193 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_62_T_2[36]}},_output_mat_62_T_2}) :
    $signed(_GEN_128); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [43:0] _GEN_194 = counter_ccnt == counter_cend ? $signed({{7{_output_mat_63_T_2[36]}},_output_mat_63_T_2}) :
    $signed(_GEN_129); // @[accumu.scala 43:46 accumu.scala 46:35]
  wire [9:0] _GEN_195 = counter_ccnt == counter_cend ? _counter_ccnt_T_1 : _GEN_65; // @[accumu.scala 43:46 accumu.scala 47:30]
  wire [43:0] _GEN_196 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_1); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_197 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_2); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_198 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_3); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_199 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_4); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_200 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_5); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_201 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_6); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_202 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_7); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_203 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_8); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_204 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_9); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_205 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_10); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_206 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_11); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_207 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_12); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_208 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_13); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_209 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_14); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_210 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_15); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_211 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_16); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_212 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_17); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_213 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_18); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_214 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_19); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_215 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_20); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_216 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_21); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_217 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_22); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_218 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_23); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_219 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_24); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_220 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_25); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_221 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_26); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_222 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_27); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_223 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_28); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_224 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_29); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_225 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_30); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_226 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_31); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_227 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_32); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_228 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_33); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_229 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_34); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_230 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_35); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_231 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_36); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_232 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_37); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_233 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_38); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_234 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_39); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_235 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_40); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_236 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_41); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_237 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_42); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_238 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_43); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_239 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_44); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_240 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_45); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_241 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_46); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_242 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_47); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_243 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_48); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_244 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_49); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_245 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_50); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_246 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_51); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_247 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_52); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_248 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_53); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_249 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_54); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_250 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_55); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_251 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_56); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_252 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_57); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_253 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_58); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_254 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_59); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_255 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_60); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_256 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_61); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_257 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_62); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_258 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_63); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire [43:0] _GEN_259 = counter_ccnt == counter_cend ? $signed(44'sh0) : $signed(_GEN_64); // @[accumu.scala 43:46 accumu.scala 32:15]
  wire  nxt = now_addr_ccnt == now_addr_cend; // @[utils.scala 17:20]
  wire [9:0] _now_addr_ccnt_T_1 = now_addr_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _now_addr_ccnt_T_2 = nxt ? 10'h0 : _now_addr_ccnt_T_1; // @[utils.scala 18:20]
  wire [9:0] _GEN_260 = counter_ccnt == 10'h1 ? _now_addr_ccnt_T_2 : now_addr_ccnt; // @[accumu.scala 59:37 utils.scala 18:14 accumu.scala 29:27]
  wire  _GEN_261 = io_valid_in & _GEN_130; // @[accumu.scala 42:26 accumu.scala 33:18]
  wire [43:0] _GEN_327 = io_valid_in ? $signed(_GEN_196) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_328 = io_valid_in ? $signed(_GEN_197) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_329 = io_valid_in ? $signed(_GEN_198) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_330 = io_valid_in ? $signed(_GEN_199) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_331 = io_valid_in ? $signed(_GEN_200) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_332 = io_valid_in ? $signed(_GEN_201) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_333 = io_valid_in ? $signed(_GEN_202) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_334 = io_valid_in ? $signed(_GEN_203) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_335 = io_valid_in ? $signed(_GEN_204) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_336 = io_valid_in ? $signed(_GEN_205) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_337 = io_valid_in ? $signed(_GEN_206) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_338 = io_valid_in ? $signed(_GEN_207) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_339 = io_valid_in ? $signed(_GEN_208) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_340 = io_valid_in ? $signed(_GEN_209) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_341 = io_valid_in ? $signed(_GEN_210) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_342 = io_valid_in ? $signed(_GEN_211) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_343 = io_valid_in ? $signed(_GEN_212) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_344 = io_valid_in ? $signed(_GEN_213) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_345 = io_valid_in ? $signed(_GEN_214) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_346 = io_valid_in ? $signed(_GEN_215) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_347 = io_valid_in ? $signed(_GEN_216) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_348 = io_valid_in ? $signed(_GEN_217) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_349 = io_valid_in ? $signed(_GEN_218) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_350 = io_valid_in ? $signed(_GEN_219) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_351 = io_valid_in ? $signed(_GEN_220) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_352 = io_valid_in ? $signed(_GEN_221) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_353 = io_valid_in ? $signed(_GEN_222) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_354 = io_valid_in ? $signed(_GEN_223) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_355 = io_valid_in ? $signed(_GEN_224) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_356 = io_valid_in ? $signed(_GEN_225) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_357 = io_valid_in ? $signed(_GEN_226) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_358 = io_valid_in ? $signed(_GEN_227) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_359 = io_valid_in ? $signed(_GEN_228) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_360 = io_valid_in ? $signed(_GEN_229) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_361 = io_valid_in ? $signed(_GEN_230) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_362 = io_valid_in ? $signed(_GEN_231) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_363 = io_valid_in ? $signed(_GEN_232) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_364 = io_valid_in ? $signed(_GEN_233) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_365 = io_valid_in ? $signed(_GEN_234) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_366 = io_valid_in ? $signed(_GEN_235) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_367 = io_valid_in ? $signed(_GEN_236) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_368 = io_valid_in ? $signed(_GEN_237) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_369 = io_valid_in ? $signed(_GEN_238) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_370 = io_valid_in ? $signed(_GEN_239) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_371 = io_valid_in ? $signed(_GEN_240) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_372 = io_valid_in ? $signed(_GEN_241) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_373 = io_valid_in ? $signed(_GEN_242) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_374 = io_valid_in ? $signed(_GEN_243) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_375 = io_valid_in ? $signed(_GEN_244) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_376 = io_valid_in ? $signed(_GEN_245) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_377 = io_valid_in ? $signed(_GEN_246) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_378 = io_valid_in ? $signed(_GEN_247) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_379 = io_valid_in ? $signed(_GEN_248) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_380 = io_valid_in ? $signed(_GEN_249) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_381 = io_valid_in ? $signed(_GEN_250) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_382 = io_valid_in ? $signed(_GEN_251) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_383 = io_valid_in ? $signed(_GEN_252) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_384 = io_valid_in ? $signed(_GEN_253) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_385 = io_valid_in ? $signed(_GEN_254) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_386 = io_valid_in ? $signed(_GEN_255) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_387 = io_valid_in ? $signed(_GEN_256) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_388 = io_valid_in ? $signed(_GEN_257) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_389 = io_valid_in ? $signed(_GEN_258) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire [43:0] _GEN_390 = io_valid_in ? $signed(_GEN_259) : $signed(44'sh0); // @[accumu.scala 42:26 accumu.scala 32:15]
  wire  _GEN_392 = enable & _GEN_261; // @[accumu.scala 41:23 accumu.scala 33:18]
  wire [43:0] _GEN_458 = enable ? $signed(_GEN_327) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_459 = enable ? $signed(_GEN_328) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_460 = enable ? $signed(_GEN_329) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_461 = enable ? $signed(_GEN_330) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_462 = enable ? $signed(_GEN_331) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_463 = enable ? $signed(_GEN_332) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_464 = enable ? $signed(_GEN_333) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_465 = enable ? $signed(_GEN_334) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_466 = enable ? $signed(_GEN_335) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_467 = enable ? $signed(_GEN_336) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_468 = enable ? $signed(_GEN_337) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_469 = enable ? $signed(_GEN_338) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_470 = enable ? $signed(_GEN_339) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_471 = enable ? $signed(_GEN_340) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_472 = enable ? $signed(_GEN_341) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_473 = enable ? $signed(_GEN_342) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_474 = enable ? $signed(_GEN_343) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_475 = enable ? $signed(_GEN_344) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_476 = enable ? $signed(_GEN_345) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_477 = enable ? $signed(_GEN_346) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_478 = enable ? $signed(_GEN_347) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_479 = enable ? $signed(_GEN_348) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_480 = enable ? $signed(_GEN_349) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_481 = enable ? $signed(_GEN_350) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_482 = enable ? $signed(_GEN_351) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_483 = enable ? $signed(_GEN_352) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_484 = enable ? $signed(_GEN_353) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_485 = enable ? $signed(_GEN_354) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_486 = enable ? $signed(_GEN_355) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_487 = enable ? $signed(_GEN_356) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_488 = enable ? $signed(_GEN_357) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_489 = enable ? $signed(_GEN_358) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_490 = enable ? $signed(_GEN_359) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_491 = enable ? $signed(_GEN_360) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_492 = enable ? $signed(_GEN_361) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_493 = enable ? $signed(_GEN_362) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_494 = enable ? $signed(_GEN_363) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_495 = enable ? $signed(_GEN_364) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_496 = enable ? $signed(_GEN_365) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_497 = enable ? $signed(_GEN_366) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_498 = enable ? $signed(_GEN_367) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_499 = enable ? $signed(_GEN_368) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_500 = enable ? $signed(_GEN_369) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_501 = enable ? $signed(_GEN_370) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_502 = enable ? $signed(_GEN_371) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_503 = enable ? $signed(_GEN_372) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_504 = enable ? $signed(_GEN_373) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_505 = enable ? $signed(_GEN_374) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_506 = enable ? $signed(_GEN_375) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_507 = enable ? $signed(_GEN_376) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_508 = enable ? $signed(_GEN_377) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_509 = enable ? $signed(_GEN_378) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_510 = enable ? $signed(_GEN_379) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_511 = enable ? $signed(_GEN_380) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_512 = enable ? $signed(_GEN_381) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_513 = enable ? $signed(_GEN_382) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_514 = enable ? $signed(_GEN_383) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_515 = enable ? $signed(_GEN_384) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_516 = enable ? $signed(_GEN_385) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_517 = enable ? $signed(_GEN_386) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_518 = enable ? $signed(_GEN_387) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_519 = enable ? $signed(_GEN_388) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_520 = enable ? $signed(_GEN_389) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  wire [43:0] _GEN_521 = enable ? $signed(_GEN_390) : $signed(44'sh0); // @[accumu.scala 41:23 accumu.scala 32:15]
  assign io_valid_out = io_flag_job ? 1'h0 : _GEN_392; // @[accumu.scala 36:22 accumu.scala 33:18]
  assign io_result_mat_0 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_458); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_1 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_459); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_2 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_460); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_3 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_461); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_4 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_462); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_5 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_463); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_6 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_464); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_7 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_465); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_8 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_466); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_9 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_467); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_10 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_468); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_11 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_469); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_12 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_470); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_13 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_471); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_14 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_472); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_15 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_473); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_16 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_474); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_17 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_475); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_18 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_476); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_19 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_477); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_20 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_478); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_21 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_479); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_22 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_480); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_23 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_481); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_24 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_482); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_25 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_483); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_26 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_484); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_27 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_485); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_28 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_486); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_29 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_487); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_30 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_488); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_31 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_489); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_32 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_490); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_33 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_491); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_34 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_492); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_35 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_493); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_36 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_494); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_37 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_495); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_38 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_496); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_39 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_497); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_40 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_498); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_41 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_499); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_42 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_500); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_43 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_501); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_44 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_502); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_45 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_503); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_46 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_504); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_47 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_505); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_48 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_506); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_49 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_507); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_50 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_508); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_51 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_509); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_52 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_510); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_53 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_511); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_54 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_512); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_55 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_513); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_56 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_514); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_57 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_515); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_58 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_516); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_59 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_517); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_60 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_518); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_61 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_519); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_62 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_520); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_result_mat_63 = io_flag_job ? $signed(44'sh0) : $signed(_GEN_521); // @[accumu.scala 36:22 accumu.scala 32:15]
  assign io_bias_addr = now_addr_ccnt; // @[accumu.scala 34:18]
  always @(posedge clock) begin
    if (reset) begin // @[accumu.scala 27:26]
      counter_ccnt <= 10'h0; // @[accumu.scala 27:26]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      counter_ccnt <= io_csum; // @[utils.scala 27:14]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        counter_ccnt <= _GEN_195;
      end
    end
    if (reset) begin // @[accumu.scala 27:26]
      counter_cend <= 10'h0; // @[accumu.scala 27:26]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      counter_cend <= io_csum; // @[utils.scala 26:14]
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_0 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_0 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_0 <= _GEN_131;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_1 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_1 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_1 <= _GEN_132;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_2 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_2 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_2 <= _GEN_133;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_3 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_3 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_3 <= _GEN_134;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_4 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_4 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_4 <= _GEN_135;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_5 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_5 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_5 <= _GEN_136;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_6 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_6 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_6 <= _GEN_137;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_7 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_7 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_7 <= _GEN_138;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_8 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_8 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_8 <= _GEN_139;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_9 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_9 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_9 <= _GEN_140;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_10 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_10 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_10 <= _GEN_141;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_11 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_11 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_11 <= _GEN_142;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_12 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_12 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_12 <= _GEN_143;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_13 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_13 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_13 <= _GEN_144;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_14 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_14 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_14 <= _GEN_145;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_15 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_15 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_15 <= _GEN_146;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_16 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_16 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_16 <= _GEN_147;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_17 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_17 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_17 <= _GEN_148;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_18 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_18 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_18 <= _GEN_149;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_19 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_19 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_19 <= _GEN_150;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_20 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_20 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_20 <= _GEN_151;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_21 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_21 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_21 <= _GEN_152;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_22 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_22 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_22 <= _GEN_153;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_23 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_23 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_23 <= _GEN_154;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_24 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_24 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_24 <= _GEN_155;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_25 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_25 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_25 <= _GEN_156;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_26 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_26 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_26 <= _GEN_157;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_27 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_27 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_27 <= _GEN_158;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_28 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_28 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_28 <= _GEN_159;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_29 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_29 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_29 <= _GEN_160;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_30 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_30 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_30 <= _GEN_161;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_31 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_31 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_31 <= _GEN_162;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_32 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_32 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_32 <= _GEN_163;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_33 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_33 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_33 <= _GEN_164;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_34 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_34 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_34 <= _GEN_165;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_35 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_35 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_35 <= _GEN_166;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_36 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_36 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_36 <= _GEN_167;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_37 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_37 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_37 <= _GEN_168;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_38 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_38 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_38 <= _GEN_169;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_39 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_39 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_39 <= _GEN_170;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_40 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_40 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_40 <= _GEN_171;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_41 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_41 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_41 <= _GEN_172;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_42 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_42 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_42 <= _GEN_173;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_43 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_43 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_43 <= _GEN_174;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_44 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_44 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_44 <= _GEN_175;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_45 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_45 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_45 <= _GEN_176;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_46 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_46 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_46 <= _GEN_177;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_47 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_47 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_47 <= _GEN_178;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_48 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_48 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_48 <= _GEN_179;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_49 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_49 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_49 <= _GEN_180;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_50 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_50 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_50 <= _GEN_181;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_51 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_51 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_51 <= _GEN_182;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_52 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_52 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_52 <= _GEN_183;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_53 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_53 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_53 <= _GEN_184;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_54 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_54 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_54 <= _GEN_185;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_55 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_55 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_55 <= _GEN_186;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_56 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_56 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_56 <= _GEN_187;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_57 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_57 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_57 <= _GEN_188;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_58 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_58 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_58 <= _GEN_189;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_59 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_59 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_59 <= _GEN_190;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_60 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_60 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_60 <= _GEN_191;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_61 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_61 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_61 <= _GEN_192;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_62 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_62 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_62 <= _GEN_193;
      end
    end
    if (reset) begin // @[accumu.scala 28:25]
      output_mat_63 <= 44'sh0; // @[accumu.scala 28:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      output_mat_63 <= 44'sh0; // @[accumu.scala 38:16]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        output_mat_63 <= _GEN_194;
      end
    end
    if (reset) begin // @[accumu.scala 29:27]
      now_addr_ccnt <= 10'h0; // @[accumu.scala 29:27]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      now_addr_ccnt <= 10'h0; // @[utils.scala 27:14]
    end else if (enable) begin // @[accumu.scala 41:23]
      if (io_valid_in) begin // @[accumu.scala 42:26]
        now_addr_ccnt <= _GEN_260;
      end
    end
    if (reset) begin // @[accumu.scala 29:27]
      now_addr_cend <= 10'h0; // @[accumu.scala 29:27]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      now_addr_cend <= io_bias_end_addr; // @[utils.scala 26:14]
    end
    if (reset) begin // @[accumu.scala 30:25]
      enable <= 1'h0; // @[accumu.scala 30:25]
    end else if (io_flag_job) begin // @[accumu.scala 36:22]
      enable <= io_is_in_use; // @[accumu.scala 40:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter_ccnt = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  counter_cend = _RAND_1[9:0];
  _RAND_2 = {2{`RANDOM}};
  output_mat_0 = _RAND_2[43:0];
  _RAND_3 = {2{`RANDOM}};
  output_mat_1 = _RAND_3[43:0];
  _RAND_4 = {2{`RANDOM}};
  output_mat_2 = _RAND_4[43:0];
  _RAND_5 = {2{`RANDOM}};
  output_mat_3 = _RAND_5[43:0];
  _RAND_6 = {2{`RANDOM}};
  output_mat_4 = _RAND_6[43:0];
  _RAND_7 = {2{`RANDOM}};
  output_mat_5 = _RAND_7[43:0];
  _RAND_8 = {2{`RANDOM}};
  output_mat_6 = _RAND_8[43:0];
  _RAND_9 = {2{`RANDOM}};
  output_mat_7 = _RAND_9[43:0];
  _RAND_10 = {2{`RANDOM}};
  output_mat_8 = _RAND_10[43:0];
  _RAND_11 = {2{`RANDOM}};
  output_mat_9 = _RAND_11[43:0];
  _RAND_12 = {2{`RANDOM}};
  output_mat_10 = _RAND_12[43:0];
  _RAND_13 = {2{`RANDOM}};
  output_mat_11 = _RAND_13[43:0];
  _RAND_14 = {2{`RANDOM}};
  output_mat_12 = _RAND_14[43:0];
  _RAND_15 = {2{`RANDOM}};
  output_mat_13 = _RAND_15[43:0];
  _RAND_16 = {2{`RANDOM}};
  output_mat_14 = _RAND_16[43:0];
  _RAND_17 = {2{`RANDOM}};
  output_mat_15 = _RAND_17[43:0];
  _RAND_18 = {2{`RANDOM}};
  output_mat_16 = _RAND_18[43:0];
  _RAND_19 = {2{`RANDOM}};
  output_mat_17 = _RAND_19[43:0];
  _RAND_20 = {2{`RANDOM}};
  output_mat_18 = _RAND_20[43:0];
  _RAND_21 = {2{`RANDOM}};
  output_mat_19 = _RAND_21[43:0];
  _RAND_22 = {2{`RANDOM}};
  output_mat_20 = _RAND_22[43:0];
  _RAND_23 = {2{`RANDOM}};
  output_mat_21 = _RAND_23[43:0];
  _RAND_24 = {2{`RANDOM}};
  output_mat_22 = _RAND_24[43:0];
  _RAND_25 = {2{`RANDOM}};
  output_mat_23 = _RAND_25[43:0];
  _RAND_26 = {2{`RANDOM}};
  output_mat_24 = _RAND_26[43:0];
  _RAND_27 = {2{`RANDOM}};
  output_mat_25 = _RAND_27[43:0];
  _RAND_28 = {2{`RANDOM}};
  output_mat_26 = _RAND_28[43:0];
  _RAND_29 = {2{`RANDOM}};
  output_mat_27 = _RAND_29[43:0];
  _RAND_30 = {2{`RANDOM}};
  output_mat_28 = _RAND_30[43:0];
  _RAND_31 = {2{`RANDOM}};
  output_mat_29 = _RAND_31[43:0];
  _RAND_32 = {2{`RANDOM}};
  output_mat_30 = _RAND_32[43:0];
  _RAND_33 = {2{`RANDOM}};
  output_mat_31 = _RAND_33[43:0];
  _RAND_34 = {2{`RANDOM}};
  output_mat_32 = _RAND_34[43:0];
  _RAND_35 = {2{`RANDOM}};
  output_mat_33 = _RAND_35[43:0];
  _RAND_36 = {2{`RANDOM}};
  output_mat_34 = _RAND_36[43:0];
  _RAND_37 = {2{`RANDOM}};
  output_mat_35 = _RAND_37[43:0];
  _RAND_38 = {2{`RANDOM}};
  output_mat_36 = _RAND_38[43:0];
  _RAND_39 = {2{`RANDOM}};
  output_mat_37 = _RAND_39[43:0];
  _RAND_40 = {2{`RANDOM}};
  output_mat_38 = _RAND_40[43:0];
  _RAND_41 = {2{`RANDOM}};
  output_mat_39 = _RAND_41[43:0];
  _RAND_42 = {2{`RANDOM}};
  output_mat_40 = _RAND_42[43:0];
  _RAND_43 = {2{`RANDOM}};
  output_mat_41 = _RAND_43[43:0];
  _RAND_44 = {2{`RANDOM}};
  output_mat_42 = _RAND_44[43:0];
  _RAND_45 = {2{`RANDOM}};
  output_mat_43 = _RAND_45[43:0];
  _RAND_46 = {2{`RANDOM}};
  output_mat_44 = _RAND_46[43:0];
  _RAND_47 = {2{`RANDOM}};
  output_mat_45 = _RAND_47[43:0];
  _RAND_48 = {2{`RANDOM}};
  output_mat_46 = _RAND_48[43:0];
  _RAND_49 = {2{`RANDOM}};
  output_mat_47 = _RAND_49[43:0];
  _RAND_50 = {2{`RANDOM}};
  output_mat_48 = _RAND_50[43:0];
  _RAND_51 = {2{`RANDOM}};
  output_mat_49 = _RAND_51[43:0];
  _RAND_52 = {2{`RANDOM}};
  output_mat_50 = _RAND_52[43:0];
  _RAND_53 = {2{`RANDOM}};
  output_mat_51 = _RAND_53[43:0];
  _RAND_54 = {2{`RANDOM}};
  output_mat_52 = _RAND_54[43:0];
  _RAND_55 = {2{`RANDOM}};
  output_mat_53 = _RAND_55[43:0];
  _RAND_56 = {2{`RANDOM}};
  output_mat_54 = _RAND_56[43:0];
  _RAND_57 = {2{`RANDOM}};
  output_mat_55 = _RAND_57[43:0];
  _RAND_58 = {2{`RANDOM}};
  output_mat_56 = _RAND_58[43:0];
  _RAND_59 = {2{`RANDOM}};
  output_mat_57 = _RAND_59[43:0];
  _RAND_60 = {2{`RANDOM}};
  output_mat_58 = _RAND_60[43:0];
  _RAND_61 = {2{`RANDOM}};
  output_mat_59 = _RAND_61[43:0];
  _RAND_62 = {2{`RANDOM}};
  output_mat_60 = _RAND_62[43:0];
  _RAND_63 = {2{`RANDOM}};
  output_mat_61 = _RAND_63[43:0];
  _RAND_64 = {2{`RANDOM}};
  output_mat_62 = _RAND_64[43:0];
  _RAND_65 = {2{`RANDOM}};
  output_mat_63 = _RAND_65[43:0];
  _RAND_66 = {1{`RANDOM}};
  now_addr_ccnt = _RAND_66[9:0];
  _RAND_67 = {1{`RANDOM}};
  now_addr_cend = _RAND_67[9:0];
  _RAND_68 = {1{`RANDOM}};
  enable = _RAND_68[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Quant(
  input         clock,
  input         reset,
  input         io_valid_in,
  output        io_valid_out,
  input         io_flag_job,
  input  [43:0] io_in_from_accumu_mat_0,
  input  [43:0] io_in_from_accumu_mat_1,
  input  [43:0] io_in_from_accumu_mat_2,
  input  [43:0] io_in_from_accumu_mat_3,
  input  [43:0] io_in_from_accumu_mat_4,
  input  [43:0] io_in_from_accumu_mat_5,
  input  [43:0] io_in_from_accumu_mat_6,
  input  [43:0] io_in_from_accumu_mat_7,
  input  [43:0] io_in_from_accumu_mat_8,
  input  [43:0] io_in_from_accumu_mat_9,
  input  [43:0] io_in_from_accumu_mat_10,
  input  [43:0] io_in_from_accumu_mat_11,
  input  [43:0] io_in_from_accumu_mat_12,
  input  [43:0] io_in_from_accumu_mat_13,
  input  [43:0] io_in_from_accumu_mat_14,
  input  [43:0] io_in_from_accumu_mat_15,
  input  [43:0] io_in_from_accumu_mat_16,
  input  [43:0] io_in_from_accumu_mat_17,
  input  [43:0] io_in_from_accumu_mat_18,
  input  [43:0] io_in_from_accumu_mat_19,
  input  [43:0] io_in_from_accumu_mat_20,
  input  [43:0] io_in_from_accumu_mat_21,
  input  [43:0] io_in_from_accumu_mat_22,
  input  [43:0] io_in_from_accumu_mat_23,
  input  [43:0] io_in_from_accumu_mat_24,
  input  [43:0] io_in_from_accumu_mat_25,
  input  [43:0] io_in_from_accumu_mat_26,
  input  [43:0] io_in_from_accumu_mat_27,
  input  [43:0] io_in_from_accumu_mat_28,
  input  [43:0] io_in_from_accumu_mat_29,
  input  [43:0] io_in_from_accumu_mat_30,
  input  [43:0] io_in_from_accumu_mat_31,
  input  [43:0] io_in_from_accumu_mat_32,
  input  [43:0] io_in_from_accumu_mat_33,
  input  [43:0] io_in_from_accumu_mat_34,
  input  [43:0] io_in_from_accumu_mat_35,
  input  [43:0] io_in_from_accumu_mat_36,
  input  [43:0] io_in_from_accumu_mat_37,
  input  [43:0] io_in_from_accumu_mat_38,
  input  [43:0] io_in_from_accumu_mat_39,
  input  [43:0] io_in_from_accumu_mat_40,
  input  [43:0] io_in_from_accumu_mat_41,
  input  [43:0] io_in_from_accumu_mat_42,
  input  [43:0] io_in_from_accumu_mat_43,
  input  [43:0] io_in_from_accumu_mat_44,
  input  [43:0] io_in_from_accumu_mat_45,
  input  [43:0] io_in_from_accumu_mat_46,
  input  [43:0] io_in_from_accumu_mat_47,
  input  [43:0] io_in_from_accumu_mat_48,
  input  [43:0] io_in_from_accumu_mat_49,
  input  [43:0] io_in_from_accumu_mat_50,
  input  [43:0] io_in_from_accumu_mat_51,
  input  [43:0] io_in_from_accumu_mat_52,
  input  [43:0] io_in_from_accumu_mat_53,
  input  [43:0] io_in_from_accumu_mat_54,
  input  [43:0] io_in_from_accumu_mat_55,
  input  [43:0] io_in_from_accumu_mat_56,
  input  [43:0] io_in_from_accumu_mat_57,
  input  [43:0] io_in_from_accumu_mat_58,
  input  [43:0] io_in_from_accumu_mat_59,
  input  [43:0] io_in_from_accumu_mat_60,
  input  [43:0] io_in_from_accumu_mat_61,
  input  [43:0] io_in_from_accumu_mat_62,
  input  [43:0] io_in_from_accumu_mat_63,
  output [15:0] io_result_mat_0,
  output [15:0] io_result_mat_1,
  output [15:0] io_result_mat_2,
  output [15:0] io_result_mat_3,
  output [15:0] io_result_mat_4,
  output [15:0] io_result_mat_5,
  output [15:0] io_result_mat_6,
  output [15:0] io_result_mat_7,
  output [15:0] io_result_mat_8,
  output [15:0] io_result_mat_9,
  output [15:0] io_result_mat_10,
  output [15:0] io_result_mat_11,
  output [15:0] io_result_mat_12,
  output [15:0] io_result_mat_13,
  output [15:0] io_result_mat_14,
  output [15:0] io_result_mat_15,
  output [15:0] io_result_mat_16,
  output [15:0] io_result_mat_17,
  output [15:0] io_result_mat_18,
  output [15:0] io_result_mat_19,
  output [15:0] io_result_mat_20,
  output [15:0] io_result_mat_21,
  output [15:0] io_result_mat_22,
  output [15:0] io_result_mat_23,
  output [15:0] io_result_mat_24,
  output [15:0] io_result_mat_25,
  output [15:0] io_result_mat_26,
  output [15:0] io_result_mat_27,
  output [15:0] io_result_mat_28,
  output [15:0] io_result_mat_29,
  output [15:0] io_result_mat_30,
  output [15:0] io_result_mat_31,
  output [15:0] io_result_mat_32,
  output [15:0] io_result_mat_33,
  output [15:0] io_result_mat_34,
  output [15:0] io_result_mat_35,
  output [15:0] io_result_mat_36,
  output [15:0] io_result_mat_37,
  output [15:0] io_result_mat_38,
  output [15:0] io_result_mat_39,
  output [15:0] io_result_mat_40,
  output [15:0] io_result_mat_41,
  output [15:0] io_result_mat_42,
  output [15:0] io_result_mat_43,
  output [15:0] io_result_mat_44,
  output [15:0] io_result_mat_45,
  output [15:0] io_result_mat_46,
  output [15:0] io_result_mat_47,
  output [15:0] io_result_mat_48,
  output [15:0] io_result_mat_49,
  output [15:0] io_result_mat_50,
  output [15:0] io_result_mat_51,
  output [15:0] io_result_mat_52,
  output [15:0] io_result_mat_53,
  output [15:0] io_result_mat_54,
  output [15:0] io_result_mat_55,
  output [15:0] io_result_mat_56,
  output [15:0] io_result_mat_57,
  output [15:0] io_result_mat_58,
  output [15:0] io_result_mat_59,
  output [15:0] io_result_mat_60,
  output [15:0] io_result_mat_61,
  output [15:0] io_result_mat_62,
  output [15:0] io_result_mat_63,
  input  [5:0]  io_quant_in_in_q,
  input  [5:0]  io_quant_in_out_q
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] quant_in_q; // @[quant.scala 77:24]
  reg [5:0] quant_out_q; // @[quant.scala 77:24]
  wire [5:0] _io_result_mat_0_T_2 = quant_out_q - quant_in_q; // @[quant.scala 63:51]
  wire [106:0] _GEN_67 = {{63{io_in_from_accumu_mat_0[43]}},io_in_from_accumu_mat_0}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_0_ret1_T = $signed(_GEN_67) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_0_ret1 = _io_result_mat_0_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_0_T_5 = $signed(io_result_mat_0_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_0_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_0_T_6 = $signed(io_result_mat_0_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_0_T_5); // @[quant.scala 53:19]
  wire [5:0] _io_result_mat_0_T_8 = quant_in_q - quant_out_q; // @[quant.scala 63:76]
  wire [43:0] _io_result_mat_0_ret1_T_1 = $signed(io_in_from_accumu_mat_0) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_0_ret1_1 = {{20{_io_result_mat_0_ret1_T_1[43]}},_io_result_mat_0_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_0_T_11 = $signed(io_result_mat_0_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_0_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_0_T_12 = $signed(io_result_mat_0_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_0_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_0_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_0_T_6) : $signed(
    _io_result_mat_0_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_69 = {{63{io_in_from_accumu_mat_1[43]}},io_in_from_accumu_mat_1}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_1_ret1_T = $signed(_GEN_69) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_1_ret1 = _io_result_mat_1_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_1_T_5 = $signed(io_result_mat_1_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_1_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_1_T_6 = $signed(io_result_mat_1_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_1_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_1_ret1_T_1 = $signed(io_in_from_accumu_mat_1) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_1_ret1_1 = {{20{_io_result_mat_1_ret1_T_1[43]}},_io_result_mat_1_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_1_T_11 = $signed(io_result_mat_1_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_1_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_1_T_12 = $signed(io_result_mat_1_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_1_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_1_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_1_T_6) : $signed(
    _io_result_mat_1_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_71 = {{63{io_in_from_accumu_mat_2[43]}},io_in_from_accumu_mat_2}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_2_ret1_T = $signed(_GEN_71) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_2_ret1 = _io_result_mat_2_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_2_T_5 = $signed(io_result_mat_2_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_2_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_2_T_6 = $signed(io_result_mat_2_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_2_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_2_ret1_T_1 = $signed(io_in_from_accumu_mat_2) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_2_ret1_1 = {{20{_io_result_mat_2_ret1_T_1[43]}},_io_result_mat_2_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_2_T_11 = $signed(io_result_mat_2_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_2_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_2_T_12 = $signed(io_result_mat_2_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_2_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_2_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_2_T_6) : $signed(
    _io_result_mat_2_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_73 = {{63{io_in_from_accumu_mat_3[43]}},io_in_from_accumu_mat_3}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_3_ret1_T = $signed(_GEN_73) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_3_ret1 = _io_result_mat_3_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_3_T_5 = $signed(io_result_mat_3_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_3_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_3_T_6 = $signed(io_result_mat_3_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_3_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_3_ret1_T_1 = $signed(io_in_from_accumu_mat_3) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_3_ret1_1 = {{20{_io_result_mat_3_ret1_T_1[43]}},_io_result_mat_3_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_3_T_11 = $signed(io_result_mat_3_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_3_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_3_T_12 = $signed(io_result_mat_3_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_3_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_3_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_3_T_6) : $signed(
    _io_result_mat_3_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_75 = {{63{io_in_from_accumu_mat_4[43]}},io_in_from_accumu_mat_4}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_4_ret1_T = $signed(_GEN_75) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_4_ret1 = _io_result_mat_4_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_4_T_5 = $signed(io_result_mat_4_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_4_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_4_T_6 = $signed(io_result_mat_4_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_4_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_4_ret1_T_1 = $signed(io_in_from_accumu_mat_4) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_4_ret1_1 = {{20{_io_result_mat_4_ret1_T_1[43]}},_io_result_mat_4_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_4_T_11 = $signed(io_result_mat_4_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_4_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_4_T_12 = $signed(io_result_mat_4_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_4_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_4_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_4_T_6) : $signed(
    _io_result_mat_4_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_77 = {{63{io_in_from_accumu_mat_5[43]}},io_in_from_accumu_mat_5}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_5_ret1_T = $signed(_GEN_77) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_5_ret1 = _io_result_mat_5_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_5_T_5 = $signed(io_result_mat_5_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_5_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_5_T_6 = $signed(io_result_mat_5_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_5_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_5_ret1_T_1 = $signed(io_in_from_accumu_mat_5) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_5_ret1_1 = {{20{_io_result_mat_5_ret1_T_1[43]}},_io_result_mat_5_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_5_T_11 = $signed(io_result_mat_5_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_5_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_5_T_12 = $signed(io_result_mat_5_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_5_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_5_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_5_T_6) : $signed(
    _io_result_mat_5_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_79 = {{63{io_in_from_accumu_mat_6[43]}},io_in_from_accumu_mat_6}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_6_ret1_T = $signed(_GEN_79) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_6_ret1 = _io_result_mat_6_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_6_T_5 = $signed(io_result_mat_6_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_6_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_6_T_6 = $signed(io_result_mat_6_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_6_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_6_ret1_T_1 = $signed(io_in_from_accumu_mat_6) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_6_ret1_1 = {{20{_io_result_mat_6_ret1_T_1[43]}},_io_result_mat_6_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_6_T_11 = $signed(io_result_mat_6_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_6_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_6_T_12 = $signed(io_result_mat_6_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_6_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_6_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_6_T_6) : $signed(
    _io_result_mat_6_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_81 = {{63{io_in_from_accumu_mat_7[43]}},io_in_from_accumu_mat_7}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_7_ret1_T = $signed(_GEN_81) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_7_ret1 = _io_result_mat_7_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_7_T_5 = $signed(io_result_mat_7_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_7_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_7_T_6 = $signed(io_result_mat_7_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_7_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_7_ret1_T_1 = $signed(io_in_from_accumu_mat_7) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_7_ret1_1 = {{20{_io_result_mat_7_ret1_T_1[43]}},_io_result_mat_7_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_7_T_11 = $signed(io_result_mat_7_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_7_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_7_T_12 = $signed(io_result_mat_7_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_7_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_7_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_7_T_6) : $signed(
    _io_result_mat_7_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_83 = {{63{io_in_from_accumu_mat_8[43]}},io_in_from_accumu_mat_8}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_8_ret1_T = $signed(_GEN_83) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_8_ret1 = _io_result_mat_8_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_8_T_5 = $signed(io_result_mat_8_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_8_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_8_T_6 = $signed(io_result_mat_8_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_8_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_8_ret1_T_1 = $signed(io_in_from_accumu_mat_8) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_8_ret1_1 = {{20{_io_result_mat_8_ret1_T_1[43]}},_io_result_mat_8_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_8_T_11 = $signed(io_result_mat_8_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_8_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_8_T_12 = $signed(io_result_mat_8_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_8_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_8_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_8_T_6) : $signed(
    _io_result_mat_8_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_85 = {{63{io_in_from_accumu_mat_9[43]}},io_in_from_accumu_mat_9}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_9_ret1_T = $signed(_GEN_85) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_9_ret1 = _io_result_mat_9_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_9_T_5 = $signed(io_result_mat_9_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_9_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_9_T_6 = $signed(io_result_mat_9_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_9_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_9_ret1_T_1 = $signed(io_in_from_accumu_mat_9) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_9_ret1_1 = {{20{_io_result_mat_9_ret1_T_1[43]}},_io_result_mat_9_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_9_T_11 = $signed(io_result_mat_9_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_9_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_9_T_12 = $signed(io_result_mat_9_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_9_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_9_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_9_T_6) : $signed(
    _io_result_mat_9_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_87 = {{63{io_in_from_accumu_mat_10[43]}},io_in_from_accumu_mat_10}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_10_ret1_T = $signed(_GEN_87) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_10_ret1 = _io_result_mat_10_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_10_T_5 = $signed(io_result_mat_10_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_10_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_10_T_6 = $signed(io_result_mat_10_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_10_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_10_ret1_T_1 = $signed(io_in_from_accumu_mat_10) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_10_ret1_1 = {{20{_io_result_mat_10_ret1_T_1[43]}},_io_result_mat_10_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_10_T_11 = $signed(io_result_mat_10_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_10_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_10_T_12 = $signed(io_result_mat_10_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_10_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_10_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_10_T_6) : $signed(
    _io_result_mat_10_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_89 = {{63{io_in_from_accumu_mat_11[43]}},io_in_from_accumu_mat_11}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_11_ret1_T = $signed(_GEN_89) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_11_ret1 = _io_result_mat_11_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_11_T_5 = $signed(io_result_mat_11_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_11_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_11_T_6 = $signed(io_result_mat_11_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_11_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_11_ret1_T_1 = $signed(io_in_from_accumu_mat_11) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_11_ret1_1 = {{20{_io_result_mat_11_ret1_T_1[43]}},_io_result_mat_11_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_11_T_11 = $signed(io_result_mat_11_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_11_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_11_T_12 = $signed(io_result_mat_11_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_11_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_11_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_11_T_6) : $signed(
    _io_result_mat_11_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_91 = {{63{io_in_from_accumu_mat_12[43]}},io_in_from_accumu_mat_12}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_12_ret1_T = $signed(_GEN_91) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_12_ret1 = _io_result_mat_12_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_12_T_5 = $signed(io_result_mat_12_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_12_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_12_T_6 = $signed(io_result_mat_12_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_12_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_12_ret1_T_1 = $signed(io_in_from_accumu_mat_12) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_12_ret1_1 = {{20{_io_result_mat_12_ret1_T_1[43]}},_io_result_mat_12_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_12_T_11 = $signed(io_result_mat_12_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_12_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_12_T_12 = $signed(io_result_mat_12_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_12_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_12_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_12_T_6) : $signed(
    _io_result_mat_12_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_93 = {{63{io_in_from_accumu_mat_13[43]}},io_in_from_accumu_mat_13}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_13_ret1_T = $signed(_GEN_93) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_13_ret1 = _io_result_mat_13_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_13_T_5 = $signed(io_result_mat_13_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_13_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_13_T_6 = $signed(io_result_mat_13_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_13_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_13_ret1_T_1 = $signed(io_in_from_accumu_mat_13) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_13_ret1_1 = {{20{_io_result_mat_13_ret1_T_1[43]}},_io_result_mat_13_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_13_T_11 = $signed(io_result_mat_13_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_13_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_13_T_12 = $signed(io_result_mat_13_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_13_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_13_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_13_T_6) : $signed(
    _io_result_mat_13_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_95 = {{63{io_in_from_accumu_mat_14[43]}},io_in_from_accumu_mat_14}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_14_ret1_T = $signed(_GEN_95) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_14_ret1 = _io_result_mat_14_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_14_T_5 = $signed(io_result_mat_14_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_14_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_14_T_6 = $signed(io_result_mat_14_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_14_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_14_ret1_T_1 = $signed(io_in_from_accumu_mat_14) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_14_ret1_1 = {{20{_io_result_mat_14_ret1_T_1[43]}},_io_result_mat_14_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_14_T_11 = $signed(io_result_mat_14_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_14_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_14_T_12 = $signed(io_result_mat_14_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_14_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_14_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_14_T_6) : $signed(
    _io_result_mat_14_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_97 = {{63{io_in_from_accumu_mat_15[43]}},io_in_from_accumu_mat_15}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_15_ret1_T = $signed(_GEN_97) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_15_ret1 = _io_result_mat_15_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_15_T_5 = $signed(io_result_mat_15_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_15_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_15_T_6 = $signed(io_result_mat_15_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_15_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_15_ret1_T_1 = $signed(io_in_from_accumu_mat_15) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_15_ret1_1 = {{20{_io_result_mat_15_ret1_T_1[43]}},_io_result_mat_15_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_15_T_11 = $signed(io_result_mat_15_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_15_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_15_T_12 = $signed(io_result_mat_15_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_15_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_15_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_15_T_6) : $signed(
    _io_result_mat_15_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_99 = {{63{io_in_from_accumu_mat_16[43]}},io_in_from_accumu_mat_16}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_16_ret1_T = $signed(_GEN_99) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_16_ret1 = _io_result_mat_16_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_16_T_5 = $signed(io_result_mat_16_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_16_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_16_T_6 = $signed(io_result_mat_16_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_16_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_16_ret1_T_1 = $signed(io_in_from_accumu_mat_16) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_16_ret1_1 = {{20{_io_result_mat_16_ret1_T_1[43]}},_io_result_mat_16_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_16_T_11 = $signed(io_result_mat_16_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_16_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_16_T_12 = $signed(io_result_mat_16_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_16_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_16_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_16_T_6) : $signed(
    _io_result_mat_16_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_101 = {{63{io_in_from_accumu_mat_17[43]}},io_in_from_accumu_mat_17}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_17_ret1_T = $signed(_GEN_101) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_17_ret1 = _io_result_mat_17_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_17_T_5 = $signed(io_result_mat_17_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_17_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_17_T_6 = $signed(io_result_mat_17_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_17_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_17_ret1_T_1 = $signed(io_in_from_accumu_mat_17) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_17_ret1_1 = {{20{_io_result_mat_17_ret1_T_1[43]}},_io_result_mat_17_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_17_T_11 = $signed(io_result_mat_17_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_17_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_17_T_12 = $signed(io_result_mat_17_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_17_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_17_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_17_T_6) : $signed(
    _io_result_mat_17_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_103 = {{63{io_in_from_accumu_mat_18[43]}},io_in_from_accumu_mat_18}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_18_ret1_T = $signed(_GEN_103) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_18_ret1 = _io_result_mat_18_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_18_T_5 = $signed(io_result_mat_18_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_18_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_18_T_6 = $signed(io_result_mat_18_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_18_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_18_ret1_T_1 = $signed(io_in_from_accumu_mat_18) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_18_ret1_1 = {{20{_io_result_mat_18_ret1_T_1[43]}},_io_result_mat_18_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_18_T_11 = $signed(io_result_mat_18_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_18_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_18_T_12 = $signed(io_result_mat_18_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_18_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_18_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_18_T_6) : $signed(
    _io_result_mat_18_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_105 = {{63{io_in_from_accumu_mat_19[43]}},io_in_from_accumu_mat_19}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_19_ret1_T = $signed(_GEN_105) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_19_ret1 = _io_result_mat_19_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_19_T_5 = $signed(io_result_mat_19_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_19_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_19_T_6 = $signed(io_result_mat_19_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_19_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_19_ret1_T_1 = $signed(io_in_from_accumu_mat_19) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_19_ret1_1 = {{20{_io_result_mat_19_ret1_T_1[43]}},_io_result_mat_19_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_19_T_11 = $signed(io_result_mat_19_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_19_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_19_T_12 = $signed(io_result_mat_19_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_19_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_19_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_19_T_6) : $signed(
    _io_result_mat_19_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_107 = {{63{io_in_from_accumu_mat_20[43]}},io_in_from_accumu_mat_20}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_20_ret1_T = $signed(_GEN_107) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_20_ret1 = _io_result_mat_20_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_20_T_5 = $signed(io_result_mat_20_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_20_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_20_T_6 = $signed(io_result_mat_20_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_20_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_20_ret1_T_1 = $signed(io_in_from_accumu_mat_20) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_20_ret1_1 = {{20{_io_result_mat_20_ret1_T_1[43]}},_io_result_mat_20_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_20_T_11 = $signed(io_result_mat_20_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_20_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_20_T_12 = $signed(io_result_mat_20_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_20_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_20_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_20_T_6) : $signed(
    _io_result_mat_20_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_109 = {{63{io_in_from_accumu_mat_21[43]}},io_in_from_accumu_mat_21}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_21_ret1_T = $signed(_GEN_109) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_21_ret1 = _io_result_mat_21_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_21_T_5 = $signed(io_result_mat_21_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_21_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_21_T_6 = $signed(io_result_mat_21_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_21_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_21_ret1_T_1 = $signed(io_in_from_accumu_mat_21) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_21_ret1_1 = {{20{_io_result_mat_21_ret1_T_1[43]}},_io_result_mat_21_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_21_T_11 = $signed(io_result_mat_21_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_21_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_21_T_12 = $signed(io_result_mat_21_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_21_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_21_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_21_T_6) : $signed(
    _io_result_mat_21_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_111 = {{63{io_in_from_accumu_mat_22[43]}},io_in_from_accumu_mat_22}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_22_ret1_T = $signed(_GEN_111) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_22_ret1 = _io_result_mat_22_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_22_T_5 = $signed(io_result_mat_22_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_22_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_22_T_6 = $signed(io_result_mat_22_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_22_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_22_ret1_T_1 = $signed(io_in_from_accumu_mat_22) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_22_ret1_1 = {{20{_io_result_mat_22_ret1_T_1[43]}},_io_result_mat_22_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_22_T_11 = $signed(io_result_mat_22_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_22_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_22_T_12 = $signed(io_result_mat_22_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_22_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_22_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_22_T_6) : $signed(
    _io_result_mat_22_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_113 = {{63{io_in_from_accumu_mat_23[43]}},io_in_from_accumu_mat_23}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_23_ret1_T = $signed(_GEN_113) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_23_ret1 = _io_result_mat_23_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_23_T_5 = $signed(io_result_mat_23_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_23_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_23_T_6 = $signed(io_result_mat_23_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_23_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_23_ret1_T_1 = $signed(io_in_from_accumu_mat_23) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_23_ret1_1 = {{20{_io_result_mat_23_ret1_T_1[43]}},_io_result_mat_23_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_23_T_11 = $signed(io_result_mat_23_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_23_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_23_T_12 = $signed(io_result_mat_23_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_23_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_23_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_23_T_6) : $signed(
    _io_result_mat_23_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_115 = {{63{io_in_from_accumu_mat_24[43]}},io_in_from_accumu_mat_24}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_24_ret1_T = $signed(_GEN_115) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_24_ret1 = _io_result_mat_24_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_24_T_5 = $signed(io_result_mat_24_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_24_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_24_T_6 = $signed(io_result_mat_24_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_24_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_24_ret1_T_1 = $signed(io_in_from_accumu_mat_24) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_24_ret1_1 = {{20{_io_result_mat_24_ret1_T_1[43]}},_io_result_mat_24_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_24_T_11 = $signed(io_result_mat_24_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_24_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_24_T_12 = $signed(io_result_mat_24_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_24_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_24_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_24_T_6) : $signed(
    _io_result_mat_24_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_117 = {{63{io_in_from_accumu_mat_25[43]}},io_in_from_accumu_mat_25}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_25_ret1_T = $signed(_GEN_117) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_25_ret1 = _io_result_mat_25_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_25_T_5 = $signed(io_result_mat_25_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_25_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_25_T_6 = $signed(io_result_mat_25_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_25_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_25_ret1_T_1 = $signed(io_in_from_accumu_mat_25) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_25_ret1_1 = {{20{_io_result_mat_25_ret1_T_1[43]}},_io_result_mat_25_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_25_T_11 = $signed(io_result_mat_25_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_25_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_25_T_12 = $signed(io_result_mat_25_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_25_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_25_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_25_T_6) : $signed(
    _io_result_mat_25_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_119 = {{63{io_in_from_accumu_mat_26[43]}},io_in_from_accumu_mat_26}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_26_ret1_T = $signed(_GEN_119) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_26_ret1 = _io_result_mat_26_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_26_T_5 = $signed(io_result_mat_26_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_26_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_26_T_6 = $signed(io_result_mat_26_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_26_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_26_ret1_T_1 = $signed(io_in_from_accumu_mat_26) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_26_ret1_1 = {{20{_io_result_mat_26_ret1_T_1[43]}},_io_result_mat_26_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_26_T_11 = $signed(io_result_mat_26_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_26_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_26_T_12 = $signed(io_result_mat_26_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_26_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_26_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_26_T_6) : $signed(
    _io_result_mat_26_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_121 = {{63{io_in_from_accumu_mat_27[43]}},io_in_from_accumu_mat_27}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_27_ret1_T = $signed(_GEN_121) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_27_ret1 = _io_result_mat_27_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_27_T_5 = $signed(io_result_mat_27_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_27_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_27_T_6 = $signed(io_result_mat_27_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_27_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_27_ret1_T_1 = $signed(io_in_from_accumu_mat_27) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_27_ret1_1 = {{20{_io_result_mat_27_ret1_T_1[43]}},_io_result_mat_27_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_27_T_11 = $signed(io_result_mat_27_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_27_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_27_T_12 = $signed(io_result_mat_27_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_27_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_27_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_27_T_6) : $signed(
    _io_result_mat_27_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_123 = {{63{io_in_from_accumu_mat_28[43]}},io_in_from_accumu_mat_28}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_28_ret1_T = $signed(_GEN_123) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_28_ret1 = _io_result_mat_28_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_28_T_5 = $signed(io_result_mat_28_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_28_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_28_T_6 = $signed(io_result_mat_28_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_28_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_28_ret1_T_1 = $signed(io_in_from_accumu_mat_28) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_28_ret1_1 = {{20{_io_result_mat_28_ret1_T_1[43]}},_io_result_mat_28_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_28_T_11 = $signed(io_result_mat_28_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_28_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_28_T_12 = $signed(io_result_mat_28_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_28_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_28_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_28_T_6) : $signed(
    _io_result_mat_28_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_125 = {{63{io_in_from_accumu_mat_29[43]}},io_in_from_accumu_mat_29}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_29_ret1_T = $signed(_GEN_125) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_29_ret1 = _io_result_mat_29_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_29_T_5 = $signed(io_result_mat_29_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_29_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_29_T_6 = $signed(io_result_mat_29_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_29_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_29_ret1_T_1 = $signed(io_in_from_accumu_mat_29) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_29_ret1_1 = {{20{_io_result_mat_29_ret1_T_1[43]}},_io_result_mat_29_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_29_T_11 = $signed(io_result_mat_29_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_29_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_29_T_12 = $signed(io_result_mat_29_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_29_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_29_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_29_T_6) : $signed(
    _io_result_mat_29_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_127 = {{63{io_in_from_accumu_mat_30[43]}},io_in_from_accumu_mat_30}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_30_ret1_T = $signed(_GEN_127) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_30_ret1 = _io_result_mat_30_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_30_T_5 = $signed(io_result_mat_30_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_30_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_30_T_6 = $signed(io_result_mat_30_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_30_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_30_ret1_T_1 = $signed(io_in_from_accumu_mat_30) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_30_ret1_1 = {{20{_io_result_mat_30_ret1_T_1[43]}},_io_result_mat_30_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_30_T_11 = $signed(io_result_mat_30_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_30_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_30_T_12 = $signed(io_result_mat_30_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_30_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_30_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_30_T_6) : $signed(
    _io_result_mat_30_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_129 = {{63{io_in_from_accumu_mat_31[43]}},io_in_from_accumu_mat_31}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_31_ret1_T = $signed(_GEN_129) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_31_ret1 = _io_result_mat_31_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_31_T_5 = $signed(io_result_mat_31_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_31_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_31_T_6 = $signed(io_result_mat_31_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_31_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_31_ret1_T_1 = $signed(io_in_from_accumu_mat_31) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_31_ret1_1 = {{20{_io_result_mat_31_ret1_T_1[43]}},_io_result_mat_31_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_31_T_11 = $signed(io_result_mat_31_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_31_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_31_T_12 = $signed(io_result_mat_31_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_31_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_31_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_31_T_6) : $signed(
    _io_result_mat_31_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_131 = {{63{io_in_from_accumu_mat_32[43]}},io_in_from_accumu_mat_32}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_32_ret1_T = $signed(_GEN_131) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_32_ret1 = _io_result_mat_32_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_32_T_5 = $signed(io_result_mat_32_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_32_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_32_T_6 = $signed(io_result_mat_32_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_32_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_32_ret1_T_1 = $signed(io_in_from_accumu_mat_32) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_32_ret1_1 = {{20{_io_result_mat_32_ret1_T_1[43]}},_io_result_mat_32_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_32_T_11 = $signed(io_result_mat_32_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_32_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_32_T_12 = $signed(io_result_mat_32_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_32_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_32_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_32_T_6) : $signed(
    _io_result_mat_32_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_133 = {{63{io_in_from_accumu_mat_33[43]}},io_in_from_accumu_mat_33}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_33_ret1_T = $signed(_GEN_133) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_33_ret1 = _io_result_mat_33_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_33_T_5 = $signed(io_result_mat_33_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_33_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_33_T_6 = $signed(io_result_mat_33_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_33_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_33_ret1_T_1 = $signed(io_in_from_accumu_mat_33) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_33_ret1_1 = {{20{_io_result_mat_33_ret1_T_1[43]}},_io_result_mat_33_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_33_T_11 = $signed(io_result_mat_33_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_33_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_33_T_12 = $signed(io_result_mat_33_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_33_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_33_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_33_T_6) : $signed(
    _io_result_mat_33_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_135 = {{63{io_in_from_accumu_mat_34[43]}},io_in_from_accumu_mat_34}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_34_ret1_T = $signed(_GEN_135) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_34_ret1 = _io_result_mat_34_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_34_T_5 = $signed(io_result_mat_34_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_34_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_34_T_6 = $signed(io_result_mat_34_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_34_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_34_ret1_T_1 = $signed(io_in_from_accumu_mat_34) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_34_ret1_1 = {{20{_io_result_mat_34_ret1_T_1[43]}},_io_result_mat_34_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_34_T_11 = $signed(io_result_mat_34_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_34_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_34_T_12 = $signed(io_result_mat_34_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_34_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_34_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_34_T_6) : $signed(
    _io_result_mat_34_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_137 = {{63{io_in_from_accumu_mat_35[43]}},io_in_from_accumu_mat_35}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_35_ret1_T = $signed(_GEN_137) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_35_ret1 = _io_result_mat_35_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_35_T_5 = $signed(io_result_mat_35_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_35_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_35_T_6 = $signed(io_result_mat_35_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_35_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_35_ret1_T_1 = $signed(io_in_from_accumu_mat_35) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_35_ret1_1 = {{20{_io_result_mat_35_ret1_T_1[43]}},_io_result_mat_35_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_35_T_11 = $signed(io_result_mat_35_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_35_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_35_T_12 = $signed(io_result_mat_35_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_35_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_35_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_35_T_6) : $signed(
    _io_result_mat_35_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_139 = {{63{io_in_from_accumu_mat_36[43]}},io_in_from_accumu_mat_36}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_36_ret1_T = $signed(_GEN_139) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_36_ret1 = _io_result_mat_36_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_36_T_5 = $signed(io_result_mat_36_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_36_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_36_T_6 = $signed(io_result_mat_36_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_36_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_36_ret1_T_1 = $signed(io_in_from_accumu_mat_36) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_36_ret1_1 = {{20{_io_result_mat_36_ret1_T_1[43]}},_io_result_mat_36_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_36_T_11 = $signed(io_result_mat_36_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_36_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_36_T_12 = $signed(io_result_mat_36_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_36_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_36_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_36_T_6) : $signed(
    _io_result_mat_36_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_141 = {{63{io_in_from_accumu_mat_37[43]}},io_in_from_accumu_mat_37}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_37_ret1_T = $signed(_GEN_141) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_37_ret1 = _io_result_mat_37_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_37_T_5 = $signed(io_result_mat_37_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_37_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_37_T_6 = $signed(io_result_mat_37_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_37_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_37_ret1_T_1 = $signed(io_in_from_accumu_mat_37) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_37_ret1_1 = {{20{_io_result_mat_37_ret1_T_1[43]}},_io_result_mat_37_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_37_T_11 = $signed(io_result_mat_37_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_37_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_37_T_12 = $signed(io_result_mat_37_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_37_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_37_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_37_T_6) : $signed(
    _io_result_mat_37_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_143 = {{63{io_in_from_accumu_mat_38[43]}},io_in_from_accumu_mat_38}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_38_ret1_T = $signed(_GEN_143) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_38_ret1 = _io_result_mat_38_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_38_T_5 = $signed(io_result_mat_38_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_38_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_38_T_6 = $signed(io_result_mat_38_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_38_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_38_ret1_T_1 = $signed(io_in_from_accumu_mat_38) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_38_ret1_1 = {{20{_io_result_mat_38_ret1_T_1[43]}},_io_result_mat_38_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_38_T_11 = $signed(io_result_mat_38_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_38_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_38_T_12 = $signed(io_result_mat_38_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_38_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_38_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_38_T_6) : $signed(
    _io_result_mat_38_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_145 = {{63{io_in_from_accumu_mat_39[43]}},io_in_from_accumu_mat_39}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_39_ret1_T = $signed(_GEN_145) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_39_ret1 = _io_result_mat_39_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_39_T_5 = $signed(io_result_mat_39_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_39_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_39_T_6 = $signed(io_result_mat_39_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_39_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_39_ret1_T_1 = $signed(io_in_from_accumu_mat_39) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_39_ret1_1 = {{20{_io_result_mat_39_ret1_T_1[43]}},_io_result_mat_39_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_39_T_11 = $signed(io_result_mat_39_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_39_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_39_T_12 = $signed(io_result_mat_39_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_39_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_39_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_39_T_6) : $signed(
    _io_result_mat_39_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_147 = {{63{io_in_from_accumu_mat_40[43]}},io_in_from_accumu_mat_40}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_40_ret1_T = $signed(_GEN_147) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_40_ret1 = _io_result_mat_40_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_40_T_5 = $signed(io_result_mat_40_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_40_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_40_T_6 = $signed(io_result_mat_40_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_40_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_40_ret1_T_1 = $signed(io_in_from_accumu_mat_40) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_40_ret1_1 = {{20{_io_result_mat_40_ret1_T_1[43]}},_io_result_mat_40_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_40_T_11 = $signed(io_result_mat_40_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_40_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_40_T_12 = $signed(io_result_mat_40_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_40_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_40_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_40_T_6) : $signed(
    _io_result_mat_40_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_149 = {{63{io_in_from_accumu_mat_41[43]}},io_in_from_accumu_mat_41}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_41_ret1_T = $signed(_GEN_149) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_41_ret1 = _io_result_mat_41_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_41_T_5 = $signed(io_result_mat_41_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_41_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_41_T_6 = $signed(io_result_mat_41_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_41_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_41_ret1_T_1 = $signed(io_in_from_accumu_mat_41) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_41_ret1_1 = {{20{_io_result_mat_41_ret1_T_1[43]}},_io_result_mat_41_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_41_T_11 = $signed(io_result_mat_41_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_41_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_41_T_12 = $signed(io_result_mat_41_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_41_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_41_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_41_T_6) : $signed(
    _io_result_mat_41_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_151 = {{63{io_in_from_accumu_mat_42[43]}},io_in_from_accumu_mat_42}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_42_ret1_T = $signed(_GEN_151) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_42_ret1 = _io_result_mat_42_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_42_T_5 = $signed(io_result_mat_42_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_42_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_42_T_6 = $signed(io_result_mat_42_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_42_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_42_ret1_T_1 = $signed(io_in_from_accumu_mat_42) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_42_ret1_1 = {{20{_io_result_mat_42_ret1_T_1[43]}},_io_result_mat_42_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_42_T_11 = $signed(io_result_mat_42_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_42_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_42_T_12 = $signed(io_result_mat_42_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_42_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_42_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_42_T_6) : $signed(
    _io_result_mat_42_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_153 = {{63{io_in_from_accumu_mat_43[43]}},io_in_from_accumu_mat_43}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_43_ret1_T = $signed(_GEN_153) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_43_ret1 = _io_result_mat_43_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_43_T_5 = $signed(io_result_mat_43_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_43_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_43_T_6 = $signed(io_result_mat_43_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_43_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_43_ret1_T_1 = $signed(io_in_from_accumu_mat_43) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_43_ret1_1 = {{20{_io_result_mat_43_ret1_T_1[43]}},_io_result_mat_43_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_43_T_11 = $signed(io_result_mat_43_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_43_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_43_T_12 = $signed(io_result_mat_43_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_43_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_43_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_43_T_6) : $signed(
    _io_result_mat_43_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_155 = {{63{io_in_from_accumu_mat_44[43]}},io_in_from_accumu_mat_44}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_44_ret1_T = $signed(_GEN_155) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_44_ret1 = _io_result_mat_44_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_44_T_5 = $signed(io_result_mat_44_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_44_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_44_T_6 = $signed(io_result_mat_44_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_44_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_44_ret1_T_1 = $signed(io_in_from_accumu_mat_44) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_44_ret1_1 = {{20{_io_result_mat_44_ret1_T_1[43]}},_io_result_mat_44_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_44_T_11 = $signed(io_result_mat_44_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_44_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_44_T_12 = $signed(io_result_mat_44_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_44_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_44_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_44_T_6) : $signed(
    _io_result_mat_44_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_157 = {{63{io_in_from_accumu_mat_45[43]}},io_in_from_accumu_mat_45}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_45_ret1_T = $signed(_GEN_157) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_45_ret1 = _io_result_mat_45_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_45_T_5 = $signed(io_result_mat_45_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_45_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_45_T_6 = $signed(io_result_mat_45_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_45_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_45_ret1_T_1 = $signed(io_in_from_accumu_mat_45) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_45_ret1_1 = {{20{_io_result_mat_45_ret1_T_1[43]}},_io_result_mat_45_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_45_T_11 = $signed(io_result_mat_45_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_45_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_45_T_12 = $signed(io_result_mat_45_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_45_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_45_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_45_T_6) : $signed(
    _io_result_mat_45_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_159 = {{63{io_in_from_accumu_mat_46[43]}},io_in_from_accumu_mat_46}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_46_ret1_T = $signed(_GEN_159) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_46_ret1 = _io_result_mat_46_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_46_T_5 = $signed(io_result_mat_46_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_46_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_46_T_6 = $signed(io_result_mat_46_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_46_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_46_ret1_T_1 = $signed(io_in_from_accumu_mat_46) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_46_ret1_1 = {{20{_io_result_mat_46_ret1_T_1[43]}},_io_result_mat_46_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_46_T_11 = $signed(io_result_mat_46_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_46_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_46_T_12 = $signed(io_result_mat_46_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_46_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_46_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_46_T_6) : $signed(
    _io_result_mat_46_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_161 = {{63{io_in_from_accumu_mat_47[43]}},io_in_from_accumu_mat_47}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_47_ret1_T = $signed(_GEN_161) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_47_ret1 = _io_result_mat_47_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_47_T_5 = $signed(io_result_mat_47_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_47_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_47_T_6 = $signed(io_result_mat_47_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_47_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_47_ret1_T_1 = $signed(io_in_from_accumu_mat_47) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_47_ret1_1 = {{20{_io_result_mat_47_ret1_T_1[43]}},_io_result_mat_47_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_47_T_11 = $signed(io_result_mat_47_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_47_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_47_T_12 = $signed(io_result_mat_47_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_47_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_47_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_47_T_6) : $signed(
    _io_result_mat_47_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_163 = {{63{io_in_from_accumu_mat_48[43]}},io_in_from_accumu_mat_48}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_48_ret1_T = $signed(_GEN_163) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_48_ret1 = _io_result_mat_48_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_48_T_5 = $signed(io_result_mat_48_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_48_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_48_T_6 = $signed(io_result_mat_48_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_48_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_48_ret1_T_1 = $signed(io_in_from_accumu_mat_48) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_48_ret1_1 = {{20{_io_result_mat_48_ret1_T_1[43]}},_io_result_mat_48_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_48_T_11 = $signed(io_result_mat_48_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_48_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_48_T_12 = $signed(io_result_mat_48_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_48_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_48_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_48_T_6) : $signed(
    _io_result_mat_48_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_165 = {{63{io_in_from_accumu_mat_49[43]}},io_in_from_accumu_mat_49}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_49_ret1_T = $signed(_GEN_165) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_49_ret1 = _io_result_mat_49_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_49_T_5 = $signed(io_result_mat_49_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_49_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_49_T_6 = $signed(io_result_mat_49_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_49_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_49_ret1_T_1 = $signed(io_in_from_accumu_mat_49) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_49_ret1_1 = {{20{_io_result_mat_49_ret1_T_1[43]}},_io_result_mat_49_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_49_T_11 = $signed(io_result_mat_49_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_49_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_49_T_12 = $signed(io_result_mat_49_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_49_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_49_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_49_T_6) : $signed(
    _io_result_mat_49_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_167 = {{63{io_in_from_accumu_mat_50[43]}},io_in_from_accumu_mat_50}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_50_ret1_T = $signed(_GEN_167) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_50_ret1 = _io_result_mat_50_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_50_T_5 = $signed(io_result_mat_50_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_50_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_50_T_6 = $signed(io_result_mat_50_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_50_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_50_ret1_T_1 = $signed(io_in_from_accumu_mat_50) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_50_ret1_1 = {{20{_io_result_mat_50_ret1_T_1[43]}},_io_result_mat_50_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_50_T_11 = $signed(io_result_mat_50_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_50_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_50_T_12 = $signed(io_result_mat_50_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_50_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_50_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_50_T_6) : $signed(
    _io_result_mat_50_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_169 = {{63{io_in_from_accumu_mat_51[43]}},io_in_from_accumu_mat_51}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_51_ret1_T = $signed(_GEN_169) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_51_ret1 = _io_result_mat_51_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_51_T_5 = $signed(io_result_mat_51_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_51_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_51_T_6 = $signed(io_result_mat_51_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_51_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_51_ret1_T_1 = $signed(io_in_from_accumu_mat_51) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_51_ret1_1 = {{20{_io_result_mat_51_ret1_T_1[43]}},_io_result_mat_51_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_51_T_11 = $signed(io_result_mat_51_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_51_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_51_T_12 = $signed(io_result_mat_51_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_51_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_51_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_51_T_6) : $signed(
    _io_result_mat_51_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_171 = {{63{io_in_from_accumu_mat_52[43]}},io_in_from_accumu_mat_52}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_52_ret1_T = $signed(_GEN_171) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_52_ret1 = _io_result_mat_52_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_52_T_5 = $signed(io_result_mat_52_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_52_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_52_T_6 = $signed(io_result_mat_52_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_52_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_52_ret1_T_1 = $signed(io_in_from_accumu_mat_52) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_52_ret1_1 = {{20{_io_result_mat_52_ret1_T_1[43]}},_io_result_mat_52_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_52_T_11 = $signed(io_result_mat_52_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_52_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_52_T_12 = $signed(io_result_mat_52_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_52_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_52_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_52_T_6) : $signed(
    _io_result_mat_52_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_173 = {{63{io_in_from_accumu_mat_53[43]}},io_in_from_accumu_mat_53}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_53_ret1_T = $signed(_GEN_173) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_53_ret1 = _io_result_mat_53_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_53_T_5 = $signed(io_result_mat_53_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_53_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_53_T_6 = $signed(io_result_mat_53_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_53_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_53_ret1_T_1 = $signed(io_in_from_accumu_mat_53) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_53_ret1_1 = {{20{_io_result_mat_53_ret1_T_1[43]}},_io_result_mat_53_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_53_T_11 = $signed(io_result_mat_53_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_53_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_53_T_12 = $signed(io_result_mat_53_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_53_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_53_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_53_T_6) : $signed(
    _io_result_mat_53_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_175 = {{63{io_in_from_accumu_mat_54[43]}},io_in_from_accumu_mat_54}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_54_ret1_T = $signed(_GEN_175) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_54_ret1 = _io_result_mat_54_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_54_T_5 = $signed(io_result_mat_54_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_54_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_54_T_6 = $signed(io_result_mat_54_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_54_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_54_ret1_T_1 = $signed(io_in_from_accumu_mat_54) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_54_ret1_1 = {{20{_io_result_mat_54_ret1_T_1[43]}},_io_result_mat_54_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_54_T_11 = $signed(io_result_mat_54_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_54_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_54_T_12 = $signed(io_result_mat_54_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_54_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_54_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_54_T_6) : $signed(
    _io_result_mat_54_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_177 = {{63{io_in_from_accumu_mat_55[43]}},io_in_from_accumu_mat_55}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_55_ret1_T = $signed(_GEN_177) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_55_ret1 = _io_result_mat_55_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_55_T_5 = $signed(io_result_mat_55_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_55_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_55_T_6 = $signed(io_result_mat_55_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_55_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_55_ret1_T_1 = $signed(io_in_from_accumu_mat_55) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_55_ret1_1 = {{20{_io_result_mat_55_ret1_T_1[43]}},_io_result_mat_55_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_55_T_11 = $signed(io_result_mat_55_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_55_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_55_T_12 = $signed(io_result_mat_55_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_55_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_55_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_55_T_6) : $signed(
    _io_result_mat_55_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_179 = {{63{io_in_from_accumu_mat_56[43]}},io_in_from_accumu_mat_56}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_56_ret1_T = $signed(_GEN_179) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_56_ret1 = _io_result_mat_56_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_56_T_5 = $signed(io_result_mat_56_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_56_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_56_T_6 = $signed(io_result_mat_56_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_56_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_56_ret1_T_1 = $signed(io_in_from_accumu_mat_56) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_56_ret1_1 = {{20{_io_result_mat_56_ret1_T_1[43]}},_io_result_mat_56_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_56_T_11 = $signed(io_result_mat_56_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_56_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_56_T_12 = $signed(io_result_mat_56_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_56_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_56_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_56_T_6) : $signed(
    _io_result_mat_56_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_181 = {{63{io_in_from_accumu_mat_57[43]}},io_in_from_accumu_mat_57}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_57_ret1_T = $signed(_GEN_181) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_57_ret1 = _io_result_mat_57_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_57_T_5 = $signed(io_result_mat_57_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_57_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_57_T_6 = $signed(io_result_mat_57_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_57_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_57_ret1_T_1 = $signed(io_in_from_accumu_mat_57) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_57_ret1_1 = {{20{_io_result_mat_57_ret1_T_1[43]}},_io_result_mat_57_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_57_T_11 = $signed(io_result_mat_57_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_57_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_57_T_12 = $signed(io_result_mat_57_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_57_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_57_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_57_T_6) : $signed(
    _io_result_mat_57_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_183 = {{63{io_in_from_accumu_mat_58[43]}},io_in_from_accumu_mat_58}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_58_ret1_T = $signed(_GEN_183) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_58_ret1 = _io_result_mat_58_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_58_T_5 = $signed(io_result_mat_58_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_58_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_58_T_6 = $signed(io_result_mat_58_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_58_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_58_ret1_T_1 = $signed(io_in_from_accumu_mat_58) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_58_ret1_1 = {{20{_io_result_mat_58_ret1_T_1[43]}},_io_result_mat_58_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_58_T_11 = $signed(io_result_mat_58_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_58_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_58_T_12 = $signed(io_result_mat_58_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_58_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_58_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_58_T_6) : $signed(
    _io_result_mat_58_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_185 = {{63{io_in_from_accumu_mat_59[43]}},io_in_from_accumu_mat_59}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_59_ret1_T = $signed(_GEN_185) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_59_ret1 = _io_result_mat_59_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_59_T_5 = $signed(io_result_mat_59_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_59_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_59_T_6 = $signed(io_result_mat_59_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_59_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_59_ret1_T_1 = $signed(io_in_from_accumu_mat_59) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_59_ret1_1 = {{20{_io_result_mat_59_ret1_T_1[43]}},_io_result_mat_59_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_59_T_11 = $signed(io_result_mat_59_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_59_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_59_T_12 = $signed(io_result_mat_59_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_59_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_59_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_59_T_6) : $signed(
    _io_result_mat_59_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_187 = {{63{io_in_from_accumu_mat_60[43]}},io_in_from_accumu_mat_60}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_60_ret1_T = $signed(_GEN_187) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_60_ret1 = _io_result_mat_60_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_60_T_5 = $signed(io_result_mat_60_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_60_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_60_T_6 = $signed(io_result_mat_60_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_60_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_60_ret1_T_1 = $signed(io_in_from_accumu_mat_60) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_60_ret1_1 = {{20{_io_result_mat_60_ret1_T_1[43]}},_io_result_mat_60_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_60_T_11 = $signed(io_result_mat_60_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_60_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_60_T_12 = $signed(io_result_mat_60_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_60_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_60_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_60_T_6) : $signed(
    _io_result_mat_60_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_189 = {{63{io_in_from_accumu_mat_61[43]}},io_in_from_accumu_mat_61}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_61_ret1_T = $signed(_GEN_189) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_61_ret1 = _io_result_mat_61_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_61_T_5 = $signed(io_result_mat_61_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_61_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_61_T_6 = $signed(io_result_mat_61_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_61_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_61_ret1_T_1 = $signed(io_in_from_accumu_mat_61) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_61_ret1_1 = {{20{_io_result_mat_61_ret1_T_1[43]}},_io_result_mat_61_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_61_T_11 = $signed(io_result_mat_61_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_61_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_61_T_12 = $signed(io_result_mat_61_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_61_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_61_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_61_T_6) : $signed(
    _io_result_mat_61_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_191 = {{63{io_in_from_accumu_mat_62[43]}},io_in_from_accumu_mat_62}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_62_ret1_T = $signed(_GEN_191) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_62_ret1 = _io_result_mat_62_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_62_T_5 = $signed(io_result_mat_62_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_62_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_62_T_6 = $signed(io_result_mat_62_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_62_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_62_ret1_T_1 = $signed(io_in_from_accumu_mat_62) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_62_ret1_1 = {{20{_io_result_mat_62_ret1_T_1[43]}},_io_result_mat_62_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_62_T_11 = $signed(io_result_mat_62_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_62_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_62_T_12 = $signed(io_result_mat_62_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_62_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_62_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_62_T_6) : $signed(
    _io_result_mat_62_T_12); // @[quant.scala 63:19]
  wire [106:0] _GEN_193 = {{63{io_in_from_accumu_mat_63[43]}},io_in_from_accumu_mat_63}; // @[quant.scala 52:18]
  wire [106:0] _io_result_mat_63_ret1_T = $signed(_GEN_193) << _io_result_mat_0_T_2; // @[quant.scala 52:18]
  wire [63:0] io_result_mat_63_ret1 = _io_result_mat_63_ret1_T[63:0]; // @[quant.scala 51:24 quant.scala 52:14]
  wire [63:0] _io_result_mat_63_T_5 = $signed(io_result_mat_63_ret1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_63_ret1); // @[quant.scala 53:41]
  wire [63:0] _io_result_mat_63_T_6 = $signed(io_result_mat_63_ret1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_63_T_5); // @[quant.scala 53:19]
  wire [43:0] _io_result_mat_63_ret1_T_1 = $signed(io_in_from_accumu_mat_63) >>> _io_result_mat_0_T_8; // @[quant.scala 59:18]
  wire [63:0] io_result_mat_63_ret1_1 = {{20{_io_result_mat_63_ret1_T_1[43]}},_io_result_mat_63_ret1_T_1}; // @[quant.scala 58:24 quant.scala 59:14]
  wire [63:0] _io_result_mat_63_T_11 = $signed(io_result_mat_63_ret1_1) >= 64'sh7fff ? $signed(64'sh7fff) : $signed(
    io_result_mat_63_ret1_1); // @[quant.scala 60:41]
  wire [63:0] _io_result_mat_63_T_12 = $signed(io_result_mat_63_ret1_1) <= -64'sh8000 ? $signed(-64'sh8000) : $signed(
    _io_result_mat_63_T_11); // @[quant.scala 60:19]
  wire [63:0] _io_result_mat_63_T_13 = quant_in_q <= quant_out_q ? $signed(_io_result_mat_63_T_6) : $signed(
    _io_result_mat_63_T_12); // @[quant.scala 63:19]
  wire [63:0] _GEN_3 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_0_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_4 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_1_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_5 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_2_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_6 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_3_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_7 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_4_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_8 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_5_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_9 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_6_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_10 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_7_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_11 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_8_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_12 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_9_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_13 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_10_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_14 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_11_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_15 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_12_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_16 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_13_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_17 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_14_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_18 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_15_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_19 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_16_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_20 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_17_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_21 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_18_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_22 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_19_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_23 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_20_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_24 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_21_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_25 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_22_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_26 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_23_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_27 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_24_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_28 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_25_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_29 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_26_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_30 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_27_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_31 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_28_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_32 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_29_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_33 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_30_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_34 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_31_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_35 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_32_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_36 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_33_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_37 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_34_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_38 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_35_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_39 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_36_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_40 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_37_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_41 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_38_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_42 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_39_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_43 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_40_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_44 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_41_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_45 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_42_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_46 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_43_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_47 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_44_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_48 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_45_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_49 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_46_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_50 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_47_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_51 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_48_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_52 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_49_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_53 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_50_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_54 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_51_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_55 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_52_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_56 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_53_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_57 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_54_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_58 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_55_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_59 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_56_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_60 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_57_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_61 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_58_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_62 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_59_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_63 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_60_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_64 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_61_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_65 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_62_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  wire [63:0] _GEN_66 = io_flag_job ? $signed(64'sh0) : $signed(_io_result_mat_63_T_13); // @[quant.scala 82:22 quant.scala 80:15 quant.scala 87:30]
  assign io_valid_out = io_flag_job ? 1'h0 : io_valid_in; // @[quant.scala 82:22 quant.scala 79:18 quant.scala 85:22]
  assign io_result_mat_0 = _GEN_3[15:0];
  assign io_result_mat_1 = _GEN_4[15:0];
  assign io_result_mat_2 = _GEN_5[15:0];
  assign io_result_mat_3 = _GEN_6[15:0];
  assign io_result_mat_4 = _GEN_7[15:0];
  assign io_result_mat_5 = _GEN_8[15:0];
  assign io_result_mat_6 = _GEN_9[15:0];
  assign io_result_mat_7 = _GEN_10[15:0];
  assign io_result_mat_8 = _GEN_11[15:0];
  assign io_result_mat_9 = _GEN_12[15:0];
  assign io_result_mat_10 = _GEN_13[15:0];
  assign io_result_mat_11 = _GEN_14[15:0];
  assign io_result_mat_12 = _GEN_15[15:0];
  assign io_result_mat_13 = _GEN_16[15:0];
  assign io_result_mat_14 = _GEN_17[15:0];
  assign io_result_mat_15 = _GEN_18[15:0];
  assign io_result_mat_16 = _GEN_19[15:0];
  assign io_result_mat_17 = _GEN_20[15:0];
  assign io_result_mat_18 = _GEN_21[15:0];
  assign io_result_mat_19 = _GEN_22[15:0];
  assign io_result_mat_20 = _GEN_23[15:0];
  assign io_result_mat_21 = _GEN_24[15:0];
  assign io_result_mat_22 = _GEN_25[15:0];
  assign io_result_mat_23 = _GEN_26[15:0];
  assign io_result_mat_24 = _GEN_27[15:0];
  assign io_result_mat_25 = _GEN_28[15:0];
  assign io_result_mat_26 = _GEN_29[15:0];
  assign io_result_mat_27 = _GEN_30[15:0];
  assign io_result_mat_28 = _GEN_31[15:0];
  assign io_result_mat_29 = _GEN_32[15:0];
  assign io_result_mat_30 = _GEN_33[15:0];
  assign io_result_mat_31 = _GEN_34[15:0];
  assign io_result_mat_32 = _GEN_35[15:0];
  assign io_result_mat_33 = _GEN_36[15:0];
  assign io_result_mat_34 = _GEN_37[15:0];
  assign io_result_mat_35 = _GEN_38[15:0];
  assign io_result_mat_36 = _GEN_39[15:0];
  assign io_result_mat_37 = _GEN_40[15:0];
  assign io_result_mat_38 = _GEN_41[15:0];
  assign io_result_mat_39 = _GEN_42[15:0];
  assign io_result_mat_40 = _GEN_43[15:0];
  assign io_result_mat_41 = _GEN_44[15:0];
  assign io_result_mat_42 = _GEN_45[15:0];
  assign io_result_mat_43 = _GEN_46[15:0];
  assign io_result_mat_44 = _GEN_47[15:0];
  assign io_result_mat_45 = _GEN_48[15:0];
  assign io_result_mat_46 = _GEN_49[15:0];
  assign io_result_mat_47 = _GEN_50[15:0];
  assign io_result_mat_48 = _GEN_51[15:0];
  assign io_result_mat_49 = _GEN_52[15:0];
  assign io_result_mat_50 = _GEN_53[15:0];
  assign io_result_mat_51 = _GEN_54[15:0];
  assign io_result_mat_52 = _GEN_55[15:0];
  assign io_result_mat_53 = _GEN_56[15:0];
  assign io_result_mat_54 = _GEN_57[15:0];
  assign io_result_mat_55 = _GEN_58[15:0];
  assign io_result_mat_56 = _GEN_59[15:0];
  assign io_result_mat_57 = _GEN_60[15:0];
  assign io_result_mat_58 = _GEN_61[15:0];
  assign io_result_mat_59 = _GEN_62[15:0];
  assign io_result_mat_60 = _GEN_63[15:0];
  assign io_result_mat_61 = _GEN_64[15:0];
  assign io_result_mat_62 = _GEN_65[15:0];
  assign io_result_mat_63 = _GEN_66[15:0];
  always @(posedge clock) begin
    if (reset) begin // @[quant.scala 77:24]
      quant_in_q <= 6'h0; // @[quant.scala 77:24]
    end else if (io_flag_job) begin // @[quant.scala 82:22]
      quant_in_q <= io_quant_in_in_q; // @[quant.scala 83:15]
    end
    if (reset) begin // @[quant.scala 77:24]
      quant_out_q <= 6'h0; // @[quant.scala 77:24]
    end else if (io_flag_job) begin // @[quant.scala 82:22]
      quant_out_q <= io_quant_in_out_q; // @[quant.scala 83:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quant_in_q = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  quant_out_q = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteSwitch(
  input         io_valid_in_0,
  output        io_valid_out,
  input  [15:0] io_input_0_mat_0,
  input  [15:0] io_input_0_mat_1,
  input  [15:0] io_input_0_mat_2,
  input  [15:0] io_input_0_mat_3,
  input  [15:0] io_input_0_mat_4,
  input  [15:0] io_input_0_mat_5,
  input  [15:0] io_input_0_mat_6,
  input  [15:0] io_input_0_mat_7,
  input  [15:0] io_input_0_mat_8,
  input  [15:0] io_input_0_mat_9,
  input  [15:0] io_input_0_mat_10,
  input  [15:0] io_input_0_mat_11,
  input  [15:0] io_input_0_mat_12,
  input  [15:0] io_input_0_mat_13,
  input  [15:0] io_input_0_mat_14,
  input  [15:0] io_input_0_mat_15,
  input  [15:0] io_input_0_mat_16,
  input  [15:0] io_input_0_mat_17,
  input  [15:0] io_input_0_mat_18,
  input  [15:0] io_input_0_mat_19,
  input  [15:0] io_input_0_mat_20,
  input  [15:0] io_input_0_mat_21,
  input  [15:0] io_input_0_mat_22,
  input  [15:0] io_input_0_mat_23,
  input  [15:0] io_input_0_mat_24,
  input  [15:0] io_input_0_mat_25,
  input  [15:0] io_input_0_mat_26,
  input  [15:0] io_input_0_mat_27,
  input  [15:0] io_input_0_mat_28,
  input  [15:0] io_input_0_mat_29,
  input  [15:0] io_input_0_mat_30,
  input  [15:0] io_input_0_mat_31,
  input  [15:0] io_input_0_mat_32,
  input  [15:0] io_input_0_mat_33,
  input  [15:0] io_input_0_mat_34,
  input  [15:0] io_input_0_mat_35,
  input  [15:0] io_input_0_mat_36,
  input  [15:0] io_input_0_mat_37,
  input  [15:0] io_input_0_mat_38,
  input  [15:0] io_input_0_mat_39,
  input  [15:0] io_input_0_mat_40,
  input  [15:0] io_input_0_mat_41,
  input  [15:0] io_input_0_mat_42,
  input  [15:0] io_input_0_mat_43,
  input  [15:0] io_input_0_mat_44,
  input  [15:0] io_input_0_mat_45,
  input  [15:0] io_input_0_mat_46,
  input  [15:0] io_input_0_mat_47,
  input  [15:0] io_input_0_mat_48,
  input  [15:0] io_input_0_mat_49,
  input  [15:0] io_input_0_mat_50,
  input  [15:0] io_input_0_mat_51,
  input  [15:0] io_input_0_mat_52,
  input  [15:0] io_input_0_mat_53,
  input  [15:0] io_input_0_mat_54,
  input  [15:0] io_input_0_mat_55,
  input  [15:0] io_input_0_mat_56,
  input  [15:0] io_input_0_mat_57,
  input  [15:0] io_input_0_mat_58,
  input  [15:0] io_input_0_mat_59,
  input  [15:0] io_input_0_mat_60,
  input  [15:0] io_input_0_mat_61,
  input  [15:0] io_input_0_mat_62,
  input  [15:0] io_input_0_mat_63,
  output [15:0] io_output_mat_0,
  output [15:0] io_output_mat_1,
  output [15:0] io_output_mat_2,
  output [15:0] io_output_mat_3,
  output [15:0] io_output_mat_4,
  output [15:0] io_output_mat_5,
  output [15:0] io_output_mat_6,
  output [15:0] io_output_mat_7,
  output [15:0] io_output_mat_8,
  output [15:0] io_output_mat_9,
  output [15:0] io_output_mat_10,
  output [15:0] io_output_mat_11,
  output [15:0] io_output_mat_12,
  output [15:0] io_output_mat_13,
  output [15:0] io_output_mat_14,
  output [15:0] io_output_mat_15,
  output [15:0] io_output_mat_16,
  output [15:0] io_output_mat_17,
  output [15:0] io_output_mat_18,
  output [15:0] io_output_mat_19,
  output [15:0] io_output_mat_20,
  output [15:0] io_output_mat_21,
  output [15:0] io_output_mat_22,
  output [15:0] io_output_mat_23,
  output [15:0] io_output_mat_24,
  output [15:0] io_output_mat_25,
  output [15:0] io_output_mat_26,
  output [15:0] io_output_mat_27,
  output [15:0] io_output_mat_28,
  output [15:0] io_output_mat_29,
  output [15:0] io_output_mat_30,
  output [15:0] io_output_mat_31,
  output [15:0] io_output_mat_32,
  output [15:0] io_output_mat_33,
  output [15:0] io_output_mat_34,
  output [15:0] io_output_mat_35,
  output [15:0] io_output_mat_36,
  output [15:0] io_output_mat_37,
  output [15:0] io_output_mat_38,
  output [15:0] io_output_mat_39,
  output [15:0] io_output_mat_40,
  output [15:0] io_output_mat_41,
  output [15:0] io_output_mat_42,
  output [15:0] io_output_mat_43,
  output [15:0] io_output_mat_44,
  output [15:0] io_output_mat_45,
  output [15:0] io_output_mat_46,
  output [15:0] io_output_mat_47,
  output [15:0] io_output_mat_48,
  output [15:0] io_output_mat_49,
  output [15:0] io_output_mat_50,
  output [15:0] io_output_mat_51,
  output [15:0] io_output_mat_52,
  output [15:0] io_output_mat_53,
  output [15:0] io_output_mat_54,
  output [15:0] io_output_mat_55,
  output [15:0] io_output_mat_56,
  output [15:0] io_output_mat_57,
  output [15:0] io_output_mat_58,
  output [15:0] io_output_mat_59,
  output [15:0] io_output_mat_60,
  output [15:0] io_output_mat_61,
  output [15:0] io_output_mat_62,
  output [15:0] io_output_mat_63
);
  assign io_valid_out = io_valid_in_0; // @[switch.scala 81:42]
  assign io_output_mat_0 = io_valid_in_0 ? $signed(io_input_0_mat_0) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_1 = io_valid_in_0 ? $signed(io_input_0_mat_1) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_2 = io_valid_in_0 ? $signed(io_input_0_mat_2) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_3 = io_valid_in_0 ? $signed(io_input_0_mat_3) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_4 = io_valid_in_0 ? $signed(io_input_0_mat_4) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_5 = io_valid_in_0 ? $signed(io_input_0_mat_5) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_6 = io_valid_in_0 ? $signed(io_input_0_mat_6) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_7 = io_valid_in_0 ? $signed(io_input_0_mat_7) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_8 = io_valid_in_0 ? $signed(io_input_0_mat_8) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_9 = io_valid_in_0 ? $signed(io_input_0_mat_9) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_10 = io_valid_in_0 ? $signed(io_input_0_mat_10) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_11 = io_valid_in_0 ? $signed(io_input_0_mat_11) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_12 = io_valid_in_0 ? $signed(io_input_0_mat_12) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_13 = io_valid_in_0 ? $signed(io_input_0_mat_13) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_14 = io_valid_in_0 ? $signed(io_input_0_mat_14) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_15 = io_valid_in_0 ? $signed(io_input_0_mat_15) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_16 = io_valid_in_0 ? $signed(io_input_0_mat_16) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_17 = io_valid_in_0 ? $signed(io_input_0_mat_17) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_18 = io_valid_in_0 ? $signed(io_input_0_mat_18) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_19 = io_valid_in_0 ? $signed(io_input_0_mat_19) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_20 = io_valid_in_0 ? $signed(io_input_0_mat_20) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_21 = io_valid_in_0 ? $signed(io_input_0_mat_21) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_22 = io_valid_in_0 ? $signed(io_input_0_mat_22) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_23 = io_valid_in_0 ? $signed(io_input_0_mat_23) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_24 = io_valid_in_0 ? $signed(io_input_0_mat_24) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_25 = io_valid_in_0 ? $signed(io_input_0_mat_25) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_26 = io_valid_in_0 ? $signed(io_input_0_mat_26) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_27 = io_valid_in_0 ? $signed(io_input_0_mat_27) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_28 = io_valid_in_0 ? $signed(io_input_0_mat_28) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_29 = io_valid_in_0 ? $signed(io_input_0_mat_29) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_30 = io_valid_in_0 ? $signed(io_input_0_mat_30) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_31 = io_valid_in_0 ? $signed(io_input_0_mat_31) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_32 = io_valid_in_0 ? $signed(io_input_0_mat_32) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_33 = io_valid_in_0 ? $signed(io_input_0_mat_33) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_34 = io_valid_in_0 ? $signed(io_input_0_mat_34) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_35 = io_valid_in_0 ? $signed(io_input_0_mat_35) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_36 = io_valid_in_0 ? $signed(io_input_0_mat_36) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_37 = io_valid_in_0 ? $signed(io_input_0_mat_37) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_38 = io_valid_in_0 ? $signed(io_input_0_mat_38) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_39 = io_valid_in_0 ? $signed(io_input_0_mat_39) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_40 = io_valid_in_0 ? $signed(io_input_0_mat_40) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_41 = io_valid_in_0 ? $signed(io_input_0_mat_41) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_42 = io_valid_in_0 ? $signed(io_input_0_mat_42) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_43 = io_valid_in_0 ? $signed(io_input_0_mat_43) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_44 = io_valid_in_0 ? $signed(io_input_0_mat_44) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_45 = io_valid_in_0 ? $signed(io_input_0_mat_45) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_46 = io_valid_in_0 ? $signed(io_input_0_mat_46) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_47 = io_valid_in_0 ? $signed(io_input_0_mat_47) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_48 = io_valid_in_0 ? $signed(io_input_0_mat_48) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_49 = io_valid_in_0 ? $signed(io_input_0_mat_49) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_50 = io_valid_in_0 ? $signed(io_input_0_mat_50) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_51 = io_valid_in_0 ? $signed(io_input_0_mat_51) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_52 = io_valid_in_0 ? $signed(io_input_0_mat_52) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_53 = io_valid_in_0 ? $signed(io_input_0_mat_53) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_54 = io_valid_in_0 ? $signed(io_input_0_mat_54) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_55 = io_valid_in_0 ? $signed(io_input_0_mat_55) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_56 = io_valid_in_0 ? $signed(io_input_0_mat_56) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_57 = io_valid_in_0 ? $signed(io_input_0_mat_57) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_58 = io_valid_in_0 ? $signed(io_input_0_mat_58) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_59 = io_valid_in_0 ? $signed(io_input_0_mat_59) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_60 = io_valid_in_0 ? $signed(io_input_0_mat_60) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_61 = io_valid_in_0 ? $signed(io_input_0_mat_61) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_62 = io_valid_in_0 ? $signed(io_input_0_mat_62) : $signed(16'sh0); // @[Mux.scala 98:16]
  assign io_output_mat_63 = io_valid_in_0 ? $signed(io_input_0_mat_63) : $signed(16'sh0); // @[Mux.scala 98:16]
endmodule
module RealWriter(
  input         clock,
  input         reset,
  input         io_valid_in,
  output        io_valid_out,
  input         io_flag_job,
  input  [15:0] io_in_from_quant_mat_0,
  input  [15:0] io_in_from_quant_mat_1,
  input  [15:0] io_in_from_quant_mat_2,
  input  [15:0] io_in_from_quant_mat_3,
  input  [15:0] io_in_from_quant_mat_4,
  input  [15:0] io_in_from_quant_mat_5,
  input  [15:0] io_in_from_quant_mat_6,
  input  [15:0] io_in_from_quant_mat_7,
  input  [15:0] io_in_from_quant_mat_8,
  input  [15:0] io_in_from_quant_mat_9,
  input  [15:0] io_in_from_quant_mat_10,
  input  [15:0] io_in_from_quant_mat_11,
  input  [15:0] io_in_from_quant_mat_12,
  input  [15:0] io_in_from_quant_mat_13,
  input  [15:0] io_in_from_quant_mat_14,
  input  [15:0] io_in_from_quant_mat_15,
  input  [15:0] io_in_from_quant_mat_16,
  input  [15:0] io_in_from_quant_mat_17,
  input  [15:0] io_in_from_quant_mat_18,
  input  [15:0] io_in_from_quant_mat_19,
  input  [15:0] io_in_from_quant_mat_20,
  input  [15:0] io_in_from_quant_mat_21,
  input  [15:0] io_in_from_quant_mat_22,
  input  [15:0] io_in_from_quant_mat_23,
  input  [15:0] io_in_from_quant_mat_24,
  input  [15:0] io_in_from_quant_mat_25,
  input  [15:0] io_in_from_quant_mat_26,
  input  [15:0] io_in_from_quant_mat_27,
  input  [15:0] io_in_from_quant_mat_28,
  input  [15:0] io_in_from_quant_mat_29,
  input  [15:0] io_in_from_quant_mat_30,
  input  [15:0] io_in_from_quant_mat_31,
  input  [15:0] io_in_from_quant_mat_32,
  input  [15:0] io_in_from_quant_mat_33,
  input  [15:0] io_in_from_quant_mat_34,
  input  [15:0] io_in_from_quant_mat_35,
  input  [15:0] io_in_from_quant_mat_36,
  input  [15:0] io_in_from_quant_mat_37,
  input  [15:0] io_in_from_quant_mat_38,
  input  [15:0] io_in_from_quant_mat_39,
  input  [15:0] io_in_from_quant_mat_40,
  input  [15:0] io_in_from_quant_mat_41,
  input  [15:0] io_in_from_quant_mat_42,
  input  [15:0] io_in_from_quant_mat_43,
  input  [15:0] io_in_from_quant_mat_44,
  input  [15:0] io_in_from_quant_mat_45,
  input  [15:0] io_in_from_quant_mat_46,
  input  [15:0] io_in_from_quant_mat_47,
  input  [15:0] io_in_from_quant_mat_48,
  input  [15:0] io_in_from_quant_mat_49,
  input  [15:0] io_in_from_quant_mat_50,
  input  [15:0] io_in_from_quant_mat_51,
  input  [15:0] io_in_from_quant_mat_52,
  input  [15:0] io_in_from_quant_mat_53,
  input  [15:0] io_in_from_quant_mat_54,
  input  [15:0] io_in_from_quant_mat_55,
  input  [15:0] io_in_from_quant_mat_56,
  input  [15:0] io_in_from_quant_mat_57,
  input  [15:0] io_in_from_quant_mat_58,
  input  [15:0] io_in_from_quant_mat_59,
  input  [15:0] io_in_from_quant_mat_60,
  input  [15:0] io_in_from_quant_mat_61,
  input  [15:0] io_in_from_quant_mat_62,
  input  [15:0] io_in_from_quant_mat_63,
  input  [9:0]  io_job_job_0_big_begin_addr,
  input  [9:0]  io_job_job_0_big_max_addr,
  input  [9:0]  io_job_job_0_big_cnt_ic_end,
  input  [9:0]  io_job_job_0_big_a,
  input  [9:0]  io_job_job_0_small_0_begin_addr,
  input  [9:0]  io_job_job_0_small_0_max_addr,
  input  [9:0]  io_job_job_0_small_0_cnt_y_end,
  input  [9:0]  io_job_job_0_small_0_cnt_ic_end,
  input  [9:0]  io_job_job_0_small_0_a,
  input  [2:0]  io_job_job_0_small_0_ano_bank_id,
  input  [9:0]  io_job_job_0_small_1_begin_addr,
  input  [9:0]  io_job_job_0_small_1_max_addr,
  input  [2:0]  io_job_job_0_small_1_bank_id,
  input  [9:0]  io_job_job_0_small_1_cnt_y_end,
  input  [9:0]  io_job_job_0_small_1_cnt_ic_end,
  input  [9:0]  io_job_job_0_small_1_a,
  input  [2:0]  io_job_job_0_small_1_ano_bank_id,
  input  [9:0]  io_job_job_1_big_begin_addr,
  input  [9:0]  io_job_job_1_big_max_addr,
  input  [2:0]  io_job_job_1_big_bank_id,
  input  [9:0]  io_job_job_1_big_cnt_ic_end,
  input  [9:0]  io_job_job_1_big_a,
  input  [9:0]  io_job_job_1_small_0_begin_addr,
  input  [9:0]  io_job_job_1_small_0_max_addr,
  input  [2:0]  io_job_job_1_small_0_bank_id,
  input  [9:0]  io_job_job_1_small_0_cnt_y_end,
  input  [9:0]  io_job_job_1_small_0_cnt_ic_end,
  input  [9:0]  io_job_job_1_small_0_a,
  input  [2:0]  io_job_job_1_small_0_ano_bank_id,
  input  [9:0]  io_job_job_1_small_1_begin_addr,
  input  [9:0]  io_job_job_1_small_1_max_addr,
  input  [2:0]  io_job_job_1_small_1_bank_id,
  input  [9:0]  io_job_job_1_small_1_cnt_y_end,
  input  [9:0]  io_job_job_1_small_1_cnt_ic_end,
  input  [9:0]  io_job_job_1_small_1_a,
  input  [2:0]  io_job_job_1_small_1_ano_bank_id,
  input  [9:0]  io_job_out_chan,
  output [15:0] io_to_bigbank_data_0,
  output [15:0] io_to_bigbank_data_1,
  output [15:0] io_to_bigbank_data_2,
  output [15:0] io_to_bigbank_data_3,
  output [15:0] io_to_bigbank_data_4,
  output [15:0] io_to_bigbank_data_5,
  output [15:0] io_to_bigbank_data_6,
  output [15:0] io_to_bigbank_data_7,
  output [15:0] io_to_bigbank_data_8,
  output [15:0] io_to_bigbank_data_9,
  output [15:0] io_to_bigbank_data_10,
  output [15:0] io_to_bigbank_data_11,
  output [15:0] io_to_bigbank_data_12,
  output [15:0] io_to_bigbank_data_13,
  output [15:0] io_to_bigbank_data_14,
  output [15:0] io_to_bigbank_data_15,
  output [15:0] io_to_bigbank_data_16,
  output [15:0] io_to_bigbank_data_17,
  output [15:0] io_to_bigbank_data_18,
  output [15:0] io_to_bigbank_data_19,
  output [15:0] io_to_bigbank_data_20,
  output [15:0] io_to_bigbank_data_21,
  output [15:0] io_to_bigbank_data_22,
  output [15:0] io_to_bigbank_data_23,
  output [15:0] io_to_bigbank_data_24,
  output [15:0] io_to_bigbank_data_25,
  output [15:0] io_to_bigbank_data_26,
  output [15:0] io_to_bigbank_data_27,
  output [15:0] io_to_bigbank_data_28,
  output [15:0] io_to_bigbank_data_29,
  output [15:0] io_to_bigbank_data_30,
  output [15:0] io_to_bigbank_data_31,
  output [15:0] io_to_bigbank_data_32,
  output [15:0] io_to_bigbank_data_33,
  output [15:0] io_to_bigbank_data_34,
  output [15:0] io_to_bigbank_data_35,
  output [15:0] io_to_bigbank_data_36,
  output [15:0] io_to_bigbank_data_37,
  output [15:0] io_to_bigbank_data_38,
  output [15:0] io_to_bigbank_data_39,
  output [15:0] io_to_bigbank_data_40,
  output [15:0] io_to_bigbank_data_41,
  output [15:0] io_to_bigbank_data_42,
  output [15:0] io_to_bigbank_data_43,
  output [15:0] io_to_bigbank_data_44,
  output [15:0] io_to_bigbank_data_45,
  output [15:0] io_to_bigbank_data_46,
  output [15:0] io_to_bigbank_data_47,
  output [15:0] io_to_smallbank_0_data_0,
  output [15:0] io_to_smallbank_0_data_1,
  output [15:0] io_to_smallbank_0_data_2,
  output [15:0] io_to_smallbank_0_data_3,
  output [15:0] io_to_smallbank_0_data_4,
  output [15:0] io_to_smallbank_0_data_5,
  output [15:0] io_to_smallbank_0_data_6,
  output [15:0] io_to_smallbank_0_data_7,
  output [15:0] io_to_smallbank_1_data_0,
  output [15:0] io_to_smallbank_1_data_1,
  output [15:0] io_to_smallbank_1_data_2,
  output [15:0] io_to_smallbank_1_data_3,
  output [15:0] io_to_smallbank_1_data_4,
  output [15:0] io_to_smallbank_1_data_5,
  output [15:0] io_to_smallbank_1_data_6,
  output [15:0] io_to_smallbank_1_data_7,
  output [9:0]  io_to_banks_addrs_0_addr,
  output [2:0]  io_to_banks_addrs_0_bank_id,
  output [9:0]  io_to_banks_addrs_1_addr,
  output [2:0]  io_to_banks_addrs_1_bank_id,
  output [9:0]  io_to_banks_addrs_2_addr,
  output [2:0]  io_to_banks_addrs_2_bank_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] gen_0_big_max_addr; // @[write.scala 71:22]
  reg [9:0] gen_0_big_now_addr; // @[write.scala 71:22]
  reg [9:0] gen_0_big_cnt_ic_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_0_big_cnt_ic_cend; // @[write.scala 71:22]
  reg [9:0] gen_0_big_a; // @[write.scala 71:22]
  reg [9:0] gen_0_small_0_max_addr; // @[write.scala 71:22]
  reg [9:0] gen_0_small_0_now_addr; // @[write.scala 71:22]
  reg [9:0] gen_0_small_0_cnt_ic_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_0_small_0_cnt_ic_cend; // @[write.scala 71:22]
  reg [9:0] gen_0_small_0_cnt_y_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_0_small_0_cnt_y_cend; // @[write.scala 71:22]
  reg [2:0] gen_0_small_0_bank_id; // @[write.scala 71:22]
  reg [9:0] gen_0_small_0_a; // @[write.scala 71:22]
  reg [2:0] gen_0_small_0_ano_bank_id; // @[write.scala 71:22]
  reg  gen_0_small_0_cnt_swap_ccnt; // @[write.scala 71:22]
  reg  gen_0_small_0_cnt_swap_cend; // @[write.scala 71:22]
  reg [9:0] gen_0_small_0_y_begin_addr; // @[write.scala 71:22]
  reg [9:0] gen_0_small_1_max_addr; // @[write.scala 71:22]
  reg [9:0] gen_0_small_1_now_addr; // @[write.scala 71:22]
  reg [9:0] gen_0_small_1_cnt_ic_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_0_small_1_cnt_ic_cend; // @[write.scala 71:22]
  reg [9:0] gen_0_small_1_cnt_y_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_0_small_1_cnt_y_cend; // @[write.scala 71:22]
  reg [2:0] gen_0_small_1_bank_id; // @[write.scala 71:22]
  reg [9:0] gen_0_small_1_a; // @[write.scala 71:22]
  reg [2:0] gen_0_small_1_ano_bank_id; // @[write.scala 71:22]
  reg  gen_0_small_1_cnt_swap_ccnt; // @[write.scala 71:22]
  reg  gen_0_small_1_cnt_swap_cend; // @[write.scala 71:22]
  reg [9:0] gen_0_small_1_y_begin_addr; // @[write.scala 71:22]
  reg [9:0] gen_1_big_max_addr; // @[write.scala 71:22]
  reg [9:0] gen_1_big_now_addr; // @[write.scala 71:22]
  reg [9:0] gen_1_big_cnt_ic_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_1_big_cnt_ic_cend; // @[write.scala 71:22]
  reg [2:0] gen_1_big_bank_id; // @[write.scala 71:22]
  reg [9:0] gen_1_big_a; // @[write.scala 71:22]
  reg [9:0] gen_1_small_0_max_addr; // @[write.scala 71:22]
  reg [9:0] gen_1_small_0_now_addr; // @[write.scala 71:22]
  reg [9:0] gen_1_small_0_cnt_ic_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_1_small_0_cnt_ic_cend; // @[write.scala 71:22]
  reg [9:0] gen_1_small_0_cnt_y_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_1_small_0_cnt_y_cend; // @[write.scala 71:22]
  reg [2:0] gen_1_small_0_bank_id; // @[write.scala 71:22]
  reg [9:0] gen_1_small_0_a; // @[write.scala 71:22]
  reg [2:0] gen_1_small_0_ano_bank_id; // @[write.scala 71:22]
  reg  gen_1_small_0_cnt_swap_ccnt; // @[write.scala 71:22]
  reg  gen_1_small_0_cnt_swap_cend; // @[write.scala 71:22]
  reg [9:0] gen_1_small_0_y_begin_addr; // @[write.scala 71:22]
  reg [9:0] gen_1_small_1_max_addr; // @[write.scala 71:22]
  reg [9:0] gen_1_small_1_now_addr; // @[write.scala 71:22]
  reg [9:0] gen_1_small_1_cnt_ic_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_1_small_1_cnt_ic_cend; // @[write.scala 71:22]
  reg [9:0] gen_1_small_1_cnt_y_ccnt; // @[write.scala 71:22]
  reg [9:0] gen_1_small_1_cnt_y_cend; // @[write.scala 71:22]
  reg [2:0] gen_1_small_1_bank_id; // @[write.scala 71:22]
  reg [9:0] gen_1_small_1_a; // @[write.scala 71:22]
  reg [2:0] gen_1_small_1_ano_bank_id; // @[write.scala 71:22]
  reg  gen_1_small_1_cnt_swap_ccnt; // @[write.scala 71:22]
  reg  gen_1_small_1_cnt_swap_cend; // @[write.scala 71:22]
  reg [9:0] gen_1_small_1_y_begin_addr; // @[write.scala 71:22]
  reg [9:0] cnt_ic_ccnt; // @[write.scala 72:25]
  reg [9:0] cnt_ic_cend; // @[write.scala 72:25]
  reg  state; // @[write.scala 73:24]
  wire [9:0] io_to_banks_ret_addrs_0_ret_addr = state ? gen_1_big_now_addr : gen_0_big_now_addr; // @[gen_addr.scala 15:18 gen_addr.scala 15:18]
  wire [9:0] io_to_banks_ret_addrs_1_ret_addr = state ? gen_1_small_0_now_addr : gen_0_small_0_now_addr; // @[gen_addr.scala 15:18 gen_addr.scala 15:18]
  wire [2:0] io_to_banks_ret_addrs_1_ret_bank_id = state ? gen_1_small_0_bank_id : gen_0_small_0_bank_id; // @[gen_addr.scala 16:21 gen_addr.scala 16:21]
  wire [9:0] io_to_banks_ret_addrs_2_ret_addr = state ? gen_1_small_1_now_addr : gen_0_small_1_now_addr; // @[gen_addr.scala 15:18 gen_addr.scala 15:18]
  wire [2:0] io_to_banks_ret_addrs_2_ret_bank_id = state ? gen_1_small_1_bank_id : gen_0_small_1_bank_id; // @[gen_addr.scala 16:21 gen_addr.scala 16:21]
  wire [9:0] _GEN_13 = state ? gen_1_big_cnt_ic_ccnt : gen_0_big_cnt_ic_ccnt; // @[utils.scala 17:20 utils.scala 17:20]
  wire [9:0] _GEN_15 = state ? gen_1_big_cnt_ic_cend : gen_0_big_cnt_ic_cend; // @[utils.scala 17:20 utils.scala 17:20]
  wire  nxt = _GEN_13 == _GEN_15; // @[utils.scala 17:20]
  wire [9:0] _gen_big_cnt_ic_ccnt_T_1 = _GEN_13 + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_big_cnt_ic_ccnt_T_2 = nxt ? 10'h0 : _gen_big_cnt_ic_ccnt_T_1; // @[utils.scala 18:20]
  wire [9:0] _GEN_19 = state ? gen_1_big_a : gen_0_big_a; // @[gen_addr.scala 284:33 gen_addr.scala 284:33]
  wire [9:0] _nxt_addr_T_1 = io_to_banks_ret_addrs_0_ret_addr + _GEN_19; // @[gen_addr.scala 284:33]
  wire [9:0] _nxt_addr_T_3 = io_to_banks_ret_addrs_0_ret_addr + 10'h1; // @[gen_addr.scala 286:33]
  wire [9:0] nxt_addr = nxt ? _nxt_addr_T_1 : _nxt_addr_T_3; // @[gen_addr.scala 283:27 gen_addr.scala 284:22 gen_addr.scala 286:22]
  wire [9:0] _GEN_22 = state ? gen_1_big_max_addr : gen_0_big_max_addr; // @[gen_addr.scala 48:18 gen_addr.scala 48:18]
  wire [9:0] _gen_big_now_addr_nxt_T_1 = nxt_addr - _GEN_22; // @[gen_addr.scala 49:24]
  wire [10:0] _gen_big_now_addr_nxt_T_2 = {{1'd0}, _gen_big_now_addr_nxt_T_1}; // @[gen_addr.scala 49:33]
  wire [9:0] gen_big_now_addr_nxt = nxt_addr >= _GEN_22 ? _gen_big_now_addr_nxt_T_2[9:0] : nxt_addr; // @[gen_addr.scala 48:29 gen_addr.scala 49:17 gen_addr.scala 51:17]
  wire [9:0] _GEN_29 = state ? gen_1_small_0_cnt_ic_ccnt : gen_0_small_0_cnt_ic_ccnt; // @[utils.scala 17:20 utils.scala 17:20]
  wire [9:0] _GEN_31 = state ? gen_1_small_0_cnt_ic_cend : gen_0_small_0_cnt_ic_cend; // @[utils.scala 17:20 utils.scala 17:20]
  wire  nxt_1 = _GEN_29 == _GEN_31; // @[utils.scala 17:20]
  wire [9:0] _gen_small_0_cnt_ic_ccnt_T_1 = _GEN_29 + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_small_0_cnt_ic_ccnt_T_2 = nxt_1 ? 10'h0 : _gen_small_0_cnt_ic_ccnt_T_1; // @[utils.scala 18:20]
  wire [9:0] _GEN_35 = state ? gen_1_small_0_cnt_y_ccnt : gen_0_small_0_cnt_y_ccnt; // @[utils.scala 17:20 utils.scala 17:20]
  wire [9:0] _GEN_37 = state ? gen_1_small_0_cnt_y_cend : gen_0_small_0_cnt_y_cend; // @[utils.scala 17:20 utils.scala 17:20]
  wire  nxt_2 = _GEN_35 == _GEN_37; // @[utils.scala 17:20]
  wire [9:0] _gen_small_0_cnt_y_ccnt_T_1 = _GEN_35 + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_small_0_cnt_y_ccnt_T_2 = nxt_2 ? 10'h0 : _gen_small_0_cnt_y_ccnt_T_1; // @[utils.scala 18:20]
  wire [9:0] _GEN_38 = ~state ? _gen_small_0_cnt_y_ccnt_T_2 : gen_0_small_0_cnt_y_ccnt; // @[utils.scala 18:14 utils.scala 18:14 write.scala 71:22]
  wire [9:0] _GEN_39 = state ? _gen_small_0_cnt_y_ccnt_T_2 : gen_1_small_0_cnt_y_ccnt; // @[utils.scala 18:14 utils.scala 18:14 write.scala 71:22]
  wire  _GEN_41 = state ? gen_1_small_0_cnt_swap_ccnt : gen_0_small_0_cnt_swap_ccnt; // @[utils.scala 17:20 utils.scala 17:20]
  wire  _GEN_43 = state ? gen_1_small_0_cnt_swap_cend : gen_0_small_0_cnt_swap_cend; // @[utils.scala 17:20 utils.scala 17:20]
  wire  nxt_3 = _GEN_41 == _GEN_43; // @[utils.scala 17:20]
  wire  _gen_small_0_cnt_swap_ccnt_T_2 = nxt_3 ? 1'h0 : _GEN_41 + 1'h1; // @[utils.scala 18:20]
  wire  _GEN_44 = ~state ? _gen_small_0_cnt_swap_ccnt_T_2 : gen_0_small_0_cnt_swap_ccnt; // @[utils.scala 18:14 utils.scala 18:14 write.scala 71:22]
  wire  _GEN_45 = state ? _gen_small_0_cnt_swap_ccnt_T_2 : gen_1_small_0_cnt_swap_ccnt; // @[utils.scala 18:14 utils.scala 18:14 write.scala 71:22]
  wire [9:0] _GEN_47 = state ? gen_1_small_0_a : gen_0_small_0_a; // @[gen_addr.scala 253:41 gen_addr.scala 253:41]
  wire [9:0] _nxt_addr_T_5 = io_to_banks_ret_addrs_1_ret_addr + _GEN_47; // @[gen_addr.scala 253:41]
  wire [9:0] _GEN_49 = state ? gen_1_small_0_max_addr : gen_0_small_0_max_addr; // @[gen_addr.scala 48:18 gen_addr.scala 48:18]
  wire [9:0] _GEN_56 = state ? gen_1_small_0_y_begin_addr : gen_0_small_0_y_begin_addr; // @[gen_addr.scala 256:30 gen_addr.scala 256:30]
  wire [9:0] _GEN_57 = nxt_3 ? _nxt_addr_T_5 : _GEN_56; // @[gen_addr.scala 252:37 gen_addr.scala 253:30 gen_addr.scala 256:30]
  wire [9:0] _GEN_68 = nxt_2 ? _GEN_57 : _nxt_addr_T_5; // @[gen_addr.scala 251:30 gen_addr.scala 261:26]
  wire [9:0] _nxt_addr_T_9 = io_to_banks_ret_addrs_1_ret_addr + 10'h1; // @[gen_addr.scala 264:33]
  wire [9:0] nxt_addr_1 = nxt_1 ? _GEN_68 : _nxt_addr_T_9; // @[gen_addr.scala 250:27 gen_addr.scala 264:22]
  wire [9:0] _gen_small_0_y_begin_addr_nxt_T_1 = nxt_addr_1 - _GEN_49; // @[gen_addr.scala 49:24]
  wire [10:0] _gen_small_0_y_begin_addr_nxt_T_2 = {{1'd0}, _gen_small_0_y_begin_addr_nxt_T_1}; // @[gen_addr.scala 49:33]
  wire [9:0] gen_small_0_y_begin_addr_nxt = nxt_addr_1 >= _GEN_49 ? _gen_small_0_y_begin_addr_nxt_T_2[9:0] : nxt_addr_1; // @[gen_addr.scala 48:29 gen_addr.scala 49:17 gen_addr.scala 51:17]
  wire [9:0] _GEN_53 = ~state ? gen_small_0_y_begin_addr_nxt : gen_0_small_0_y_begin_addr; // @[gen_addr.scala 254:34 gen_addr.scala 254:34 write.scala 71:22]
  wire [9:0] _GEN_54 = state ? gen_small_0_y_begin_addr_nxt : gen_1_small_0_y_begin_addr; // @[gen_addr.scala 254:34 gen_addr.scala 254:34 write.scala 71:22]
  wire [9:0] _GEN_58 = nxt_3 ? _GEN_53 : gen_0_small_0_y_begin_addr; // @[gen_addr.scala 252:37 write.scala 71:22]
  wire [9:0] _GEN_59 = nxt_3 ? _GEN_54 : gen_1_small_0_y_begin_addr; // @[gen_addr.scala 252:37 write.scala 71:22]
  wire [2:0] _GEN_63 = state ? gen_1_small_0_ano_bank_id : gen_0_small_0_ano_bank_id; // @[gen_addr.scala 258:25 gen_addr.scala 258:25]
  wire [2:0] _GEN_60 = ~state ? _GEN_63 : gen_0_small_0_bank_id; // @[gen_addr.scala 258:25 gen_addr.scala 258:25 write.scala 71:22]
  wire [2:0] _GEN_61 = state ? _GEN_63 : gen_1_small_0_bank_id; // @[gen_addr.scala 258:25 gen_addr.scala 258:25 write.scala 71:22]
  wire [2:0] _GEN_64 = ~state ? io_to_banks_ret_addrs_1_ret_bank_id : gen_0_small_0_ano_bank_id; // @[gen_addr.scala 259:29 gen_addr.scala 259:29 write.scala 71:22]
  wire [2:0] _GEN_65 = state ? io_to_banks_ret_addrs_1_ret_bank_id : gen_1_small_0_ano_bank_id; // @[gen_addr.scala 259:29 gen_addr.scala 259:29 write.scala 71:22]
  wire  _GEN_66 = nxt_2 ? _GEN_44 : gen_0_small_0_cnt_swap_ccnt; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire  _GEN_67 = nxt_2 ? _GEN_45 : gen_1_small_0_cnt_swap_ccnt; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [9:0] _GEN_69 = nxt_2 ? _GEN_58 : gen_0_small_0_y_begin_addr; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [9:0] _GEN_70 = nxt_2 ? _GEN_59 : gen_1_small_0_y_begin_addr; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [2:0] _GEN_71 = nxt_2 ? _GEN_60 : gen_0_small_0_bank_id; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [2:0] _GEN_72 = nxt_2 ? _GEN_61 : gen_1_small_0_bank_id; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [2:0] _GEN_73 = nxt_2 ? _GEN_64 : gen_0_small_0_ano_bank_id; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [2:0] _GEN_74 = nxt_2 ? _GEN_65 : gen_1_small_0_ano_bank_id; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [9:0] _GEN_90 = state ? gen_1_small_1_cnt_ic_ccnt : gen_0_small_1_cnt_ic_ccnt; // @[utils.scala 17:20 utils.scala 17:20]
  wire [9:0] _GEN_92 = state ? gen_1_small_1_cnt_ic_cend : gen_0_small_1_cnt_ic_cend; // @[utils.scala 17:20 utils.scala 17:20]
  wire  nxt_4 = _GEN_90 == _GEN_92; // @[utils.scala 17:20]
  wire [9:0] _gen_small_1_cnt_ic_ccnt_T_1 = _GEN_90 + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_small_1_cnt_ic_ccnt_T_2 = nxt_4 ? 10'h0 : _gen_small_1_cnt_ic_ccnt_T_1; // @[utils.scala 18:20]
  wire [9:0] _GEN_96 = state ? gen_1_small_1_cnt_y_ccnt : gen_0_small_1_cnt_y_ccnt; // @[utils.scala 17:20 utils.scala 17:20]
  wire [9:0] _GEN_98 = state ? gen_1_small_1_cnt_y_cend : gen_0_small_1_cnt_y_cend; // @[utils.scala 17:20 utils.scala 17:20]
  wire  nxt_5 = _GEN_96 == _GEN_98; // @[utils.scala 17:20]
  wire [9:0] _gen_small_1_cnt_y_ccnt_T_1 = _GEN_96 + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _gen_small_1_cnt_y_ccnt_T_2 = nxt_5 ? 10'h0 : _gen_small_1_cnt_y_ccnt_T_1; // @[utils.scala 18:20]
  wire [9:0] _GEN_99 = ~state ? _gen_small_1_cnt_y_ccnt_T_2 : gen_0_small_1_cnt_y_ccnt; // @[utils.scala 18:14 utils.scala 18:14 write.scala 71:22]
  wire [9:0] _GEN_100 = state ? _gen_small_1_cnt_y_ccnt_T_2 : gen_1_small_1_cnt_y_ccnt; // @[utils.scala 18:14 utils.scala 18:14 write.scala 71:22]
  wire  _GEN_102 = state ? gen_1_small_1_cnt_swap_ccnt : gen_0_small_1_cnt_swap_ccnt; // @[utils.scala 17:20 utils.scala 17:20]
  wire  _GEN_104 = state ? gen_1_small_1_cnt_swap_cend : gen_0_small_1_cnt_swap_cend; // @[utils.scala 17:20 utils.scala 17:20]
  wire  nxt_6 = _GEN_102 == _GEN_104; // @[utils.scala 17:20]
  wire  _gen_small_1_cnt_swap_ccnt_T_2 = nxt_6 ? 1'h0 : _GEN_102 + 1'h1; // @[utils.scala 18:20]
  wire  _GEN_105 = ~state ? _gen_small_1_cnt_swap_ccnt_T_2 : gen_0_small_1_cnt_swap_ccnt; // @[utils.scala 18:14 utils.scala 18:14 write.scala 71:22]
  wire  _GEN_106 = state ? _gen_small_1_cnt_swap_ccnt_T_2 : gen_1_small_1_cnt_swap_ccnt; // @[utils.scala 18:14 utils.scala 18:14 write.scala 71:22]
  wire [9:0] _GEN_108 = state ? gen_1_small_1_a : gen_0_small_1_a; // @[gen_addr.scala 253:41 gen_addr.scala 253:41]
  wire [9:0] _nxt_addr_T_11 = io_to_banks_ret_addrs_2_ret_addr + _GEN_108; // @[gen_addr.scala 253:41]
  wire [9:0] _GEN_110 = state ? gen_1_small_1_max_addr : gen_0_small_1_max_addr; // @[gen_addr.scala 48:18 gen_addr.scala 48:18]
  wire [9:0] _GEN_117 = state ? gen_1_small_1_y_begin_addr : gen_0_small_1_y_begin_addr; // @[gen_addr.scala 256:30 gen_addr.scala 256:30]
  wire [9:0] _GEN_118 = nxt_6 ? _nxt_addr_T_11 : _GEN_117; // @[gen_addr.scala 252:37 gen_addr.scala 253:30 gen_addr.scala 256:30]
  wire [9:0] _GEN_129 = nxt_5 ? _GEN_118 : _nxt_addr_T_11; // @[gen_addr.scala 251:30 gen_addr.scala 261:26]
  wire [9:0] _nxt_addr_T_15 = io_to_banks_ret_addrs_2_ret_addr + 10'h1; // @[gen_addr.scala 264:33]
  wire [9:0] nxt_addr_2 = nxt_4 ? _GEN_129 : _nxt_addr_T_15; // @[gen_addr.scala 250:27 gen_addr.scala 264:22]
  wire [9:0] _gen_small_1_y_begin_addr_nxt_T_1 = nxt_addr_2 - _GEN_110; // @[gen_addr.scala 49:24]
  wire [10:0] _gen_small_1_y_begin_addr_nxt_T_2 = {{1'd0}, _gen_small_1_y_begin_addr_nxt_T_1}; // @[gen_addr.scala 49:33]
  wire [9:0] gen_small_1_y_begin_addr_nxt = nxt_addr_2 >= _GEN_110 ? _gen_small_1_y_begin_addr_nxt_T_2[9:0] : nxt_addr_2
    ; // @[gen_addr.scala 48:29 gen_addr.scala 49:17 gen_addr.scala 51:17]
  wire [9:0] _GEN_114 = ~state ? gen_small_1_y_begin_addr_nxt : gen_0_small_1_y_begin_addr; // @[gen_addr.scala 254:34 gen_addr.scala 254:34 write.scala 71:22]
  wire [9:0] _GEN_115 = state ? gen_small_1_y_begin_addr_nxt : gen_1_small_1_y_begin_addr; // @[gen_addr.scala 254:34 gen_addr.scala 254:34 write.scala 71:22]
  wire [9:0] _GEN_119 = nxt_6 ? _GEN_114 : gen_0_small_1_y_begin_addr; // @[gen_addr.scala 252:37 write.scala 71:22]
  wire [9:0] _GEN_120 = nxt_6 ? _GEN_115 : gen_1_small_1_y_begin_addr; // @[gen_addr.scala 252:37 write.scala 71:22]
  wire [2:0] _GEN_124 = state ? gen_1_small_1_ano_bank_id : gen_0_small_1_ano_bank_id; // @[gen_addr.scala 258:25 gen_addr.scala 258:25]
  wire [2:0] _GEN_121 = ~state ? _GEN_124 : gen_0_small_1_bank_id; // @[gen_addr.scala 258:25 gen_addr.scala 258:25 write.scala 71:22]
  wire [2:0] _GEN_122 = state ? _GEN_124 : gen_1_small_1_bank_id; // @[gen_addr.scala 258:25 gen_addr.scala 258:25 write.scala 71:22]
  wire [2:0] _GEN_125 = ~state ? io_to_banks_ret_addrs_2_ret_bank_id : gen_0_small_1_ano_bank_id; // @[gen_addr.scala 259:29 gen_addr.scala 259:29 write.scala 71:22]
  wire [2:0] _GEN_126 = state ? io_to_banks_ret_addrs_2_ret_bank_id : gen_1_small_1_ano_bank_id; // @[gen_addr.scala 259:29 gen_addr.scala 259:29 write.scala 71:22]
  wire  _GEN_127 = nxt_5 ? _GEN_105 : gen_0_small_1_cnt_swap_ccnt; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire  _GEN_128 = nxt_5 ? _GEN_106 : gen_1_small_1_cnt_swap_ccnt; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [9:0] _GEN_130 = nxt_5 ? _GEN_119 : gen_0_small_1_y_begin_addr; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [9:0] _GEN_131 = nxt_5 ? _GEN_120 : gen_1_small_1_y_begin_addr; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [2:0] _GEN_132 = nxt_5 ? _GEN_121 : gen_0_small_1_bank_id; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [2:0] _GEN_133 = nxt_5 ? _GEN_122 : gen_1_small_1_bank_id; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [2:0] _GEN_134 = nxt_5 ? _GEN_125 : gen_0_small_1_ano_bank_id; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire [2:0] _GEN_135 = nxt_5 ? _GEN_126 : gen_1_small_1_ano_bank_id; // @[gen_addr.scala 251:30 write.scala 71:22]
  wire  nxt_7 = cnt_ic_ccnt == cnt_ic_cend; // @[utils.scala 17:20]
  wire [9:0] _cnt_ic_ccnt_T_1 = cnt_ic_ccnt + 10'h1; // @[utils.scala 18:35]
  wire  _GEN_214 = io_flag_job | gen_0_small_0_cnt_swap_cend; // @[write.scala 85:22 utils.scala 22:14 write.scala 71:22]
  wire  _GEN_231 = io_flag_job | gen_0_small_1_cnt_swap_cend; // @[write.scala 85:22 utils.scala 22:14 write.scala 71:22]
  wire  _GEN_261 = io_flag_job | gen_1_small_0_cnt_swap_cend; // @[write.scala 85:22 utils.scala 22:14 write.scala 71:22]
  wire  _GEN_278 = io_flag_job | gen_1_small_1_cnt_swap_cend; // @[write.scala 85:22 utils.scala 22:14 write.scala 71:22]
  assign io_valid_out = io_flag_job ? 1'h0 : io_valid_in; // @[write.scala 85:22 write.scala 84:18]
  assign io_to_bigbank_data_0 = io_in_from_quant_mat_1; // @[write.scala 77:39]
  assign io_to_bigbank_data_1 = io_in_from_quant_mat_2; // @[write.scala 77:39]
  assign io_to_bigbank_data_2 = io_in_from_quant_mat_3; // @[write.scala 77:39]
  assign io_to_bigbank_data_3 = io_in_from_quant_mat_4; // @[write.scala 77:39]
  assign io_to_bigbank_data_4 = io_in_from_quant_mat_5; // @[write.scala 77:39]
  assign io_to_bigbank_data_5 = io_in_from_quant_mat_6; // @[write.scala 77:39]
  assign io_to_bigbank_data_6 = io_in_from_quant_mat_9; // @[write.scala 77:39]
  assign io_to_bigbank_data_7 = io_in_from_quant_mat_10; // @[write.scala 77:39]
  assign io_to_bigbank_data_8 = io_in_from_quant_mat_11; // @[write.scala 77:39]
  assign io_to_bigbank_data_9 = io_in_from_quant_mat_12; // @[write.scala 77:39]
  assign io_to_bigbank_data_10 = io_in_from_quant_mat_13; // @[write.scala 77:39]
  assign io_to_bigbank_data_11 = io_in_from_quant_mat_14; // @[write.scala 77:39]
  assign io_to_bigbank_data_12 = io_in_from_quant_mat_17; // @[write.scala 77:39]
  assign io_to_bigbank_data_13 = io_in_from_quant_mat_18; // @[write.scala 77:39]
  assign io_to_bigbank_data_14 = io_in_from_quant_mat_19; // @[write.scala 77:39]
  assign io_to_bigbank_data_15 = io_in_from_quant_mat_20; // @[write.scala 77:39]
  assign io_to_bigbank_data_16 = io_in_from_quant_mat_21; // @[write.scala 77:39]
  assign io_to_bigbank_data_17 = io_in_from_quant_mat_22; // @[write.scala 77:39]
  assign io_to_bigbank_data_18 = io_in_from_quant_mat_25; // @[write.scala 77:39]
  assign io_to_bigbank_data_19 = io_in_from_quant_mat_26; // @[write.scala 77:39]
  assign io_to_bigbank_data_20 = io_in_from_quant_mat_27; // @[write.scala 77:39]
  assign io_to_bigbank_data_21 = io_in_from_quant_mat_28; // @[write.scala 77:39]
  assign io_to_bigbank_data_22 = io_in_from_quant_mat_29; // @[write.scala 77:39]
  assign io_to_bigbank_data_23 = io_in_from_quant_mat_30; // @[write.scala 77:39]
  assign io_to_bigbank_data_24 = io_in_from_quant_mat_33; // @[write.scala 77:39]
  assign io_to_bigbank_data_25 = io_in_from_quant_mat_34; // @[write.scala 77:39]
  assign io_to_bigbank_data_26 = io_in_from_quant_mat_35; // @[write.scala 77:39]
  assign io_to_bigbank_data_27 = io_in_from_quant_mat_36; // @[write.scala 77:39]
  assign io_to_bigbank_data_28 = io_in_from_quant_mat_37; // @[write.scala 77:39]
  assign io_to_bigbank_data_29 = io_in_from_quant_mat_38; // @[write.scala 77:39]
  assign io_to_bigbank_data_30 = io_in_from_quant_mat_41; // @[write.scala 77:39]
  assign io_to_bigbank_data_31 = io_in_from_quant_mat_42; // @[write.scala 77:39]
  assign io_to_bigbank_data_32 = io_in_from_quant_mat_43; // @[write.scala 77:39]
  assign io_to_bigbank_data_33 = io_in_from_quant_mat_44; // @[write.scala 77:39]
  assign io_to_bigbank_data_34 = io_in_from_quant_mat_45; // @[write.scala 77:39]
  assign io_to_bigbank_data_35 = io_in_from_quant_mat_46; // @[write.scala 77:39]
  assign io_to_bigbank_data_36 = io_in_from_quant_mat_49; // @[write.scala 77:39]
  assign io_to_bigbank_data_37 = io_in_from_quant_mat_50; // @[write.scala 77:39]
  assign io_to_bigbank_data_38 = io_in_from_quant_mat_51; // @[write.scala 77:39]
  assign io_to_bigbank_data_39 = io_in_from_quant_mat_52; // @[write.scala 77:39]
  assign io_to_bigbank_data_40 = io_in_from_quant_mat_53; // @[write.scala 77:39]
  assign io_to_bigbank_data_41 = io_in_from_quant_mat_54; // @[write.scala 77:39]
  assign io_to_bigbank_data_42 = io_in_from_quant_mat_57; // @[write.scala 77:39]
  assign io_to_bigbank_data_43 = io_in_from_quant_mat_58; // @[write.scala 77:39]
  assign io_to_bigbank_data_44 = io_in_from_quant_mat_59; // @[write.scala 77:39]
  assign io_to_bigbank_data_45 = io_in_from_quant_mat_60; // @[write.scala 77:39]
  assign io_to_bigbank_data_46 = io_in_from_quant_mat_61; // @[write.scala 77:39]
  assign io_to_bigbank_data_47 = io_in_from_quant_mat_62; // @[write.scala 77:39]
  assign io_to_smallbank_0_data_0 = io_in_from_quant_mat_0; // @[write.scala 79:36]
  assign io_to_smallbank_0_data_1 = io_in_from_quant_mat_8; // @[write.scala 79:36]
  assign io_to_smallbank_0_data_2 = io_in_from_quant_mat_16; // @[write.scala 79:36]
  assign io_to_smallbank_0_data_3 = io_in_from_quant_mat_24; // @[write.scala 79:36]
  assign io_to_smallbank_0_data_4 = io_in_from_quant_mat_32; // @[write.scala 79:36]
  assign io_to_smallbank_0_data_5 = io_in_from_quant_mat_40; // @[write.scala 79:36]
  assign io_to_smallbank_0_data_6 = io_in_from_quant_mat_48; // @[write.scala 79:36]
  assign io_to_smallbank_0_data_7 = io_in_from_quant_mat_56; // @[write.scala 79:36]
  assign io_to_smallbank_1_data_0 = io_in_from_quant_mat_7; // @[write.scala 81:36]
  assign io_to_smallbank_1_data_1 = io_in_from_quant_mat_15; // @[write.scala 81:36]
  assign io_to_smallbank_1_data_2 = io_in_from_quant_mat_23; // @[write.scala 81:36]
  assign io_to_smallbank_1_data_3 = io_in_from_quant_mat_31; // @[write.scala 81:36]
  assign io_to_smallbank_1_data_4 = io_in_from_quant_mat_39; // @[write.scala 81:36]
  assign io_to_smallbank_1_data_5 = io_in_from_quant_mat_47; // @[write.scala 81:36]
  assign io_to_smallbank_1_data_6 = io_in_from_quant_mat_55; // @[write.scala 81:36]
  assign io_to_smallbank_1_data_7 = io_in_from_quant_mat_63; // @[write.scala 81:36]
  assign io_to_banks_addrs_0_addr = state ? gen_1_big_now_addr : gen_0_big_now_addr; // @[gen_addr.scala 15:18 gen_addr.scala 15:18]
  assign io_to_banks_addrs_0_bank_id = state ? gen_1_big_bank_id : 3'h0; // @[gen_addr.scala 16:21 gen_addr.scala 16:21]
  assign io_to_banks_addrs_1_addr = state ? gen_1_small_0_now_addr : gen_0_small_0_now_addr; // @[gen_addr.scala 15:18 gen_addr.scala 15:18]
  assign io_to_banks_addrs_1_bank_id = state ? gen_1_small_0_bank_id : gen_0_small_0_bank_id; // @[gen_addr.scala 16:21 gen_addr.scala 16:21]
  assign io_to_banks_addrs_2_addr = state ? gen_1_small_1_now_addr : gen_0_small_1_now_addr; // @[gen_addr.scala 15:18 gen_addr.scala 15:18]
  assign io_to_banks_addrs_2_bank_id = state ? gen_1_small_1_bank_id : gen_0_small_1_bank_id; // @[gen_addr.scala 16:21 gen_addr.scala 16:21]
  always @(posedge clock) begin
    if (reset) begin // @[write.scala 71:22]
      gen_0_big_max_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_big_max_addr <= io_job_job_0_big_max_addr; // @[gen_addr.scala 56:18]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_big_now_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_big_now_addr <= io_job_job_0_big_begin_addr; // @[gen_addr.scala 58:18]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (~state) begin // @[gen_addr.scala 288:18]
        gen_0_big_now_addr <= gen_big_now_addr_nxt; // @[gen_addr.scala 288:18]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_big_cnt_ic_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_big_cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (~state) begin // @[utils.scala 18:14]
        gen_0_big_cnt_ic_ccnt <= _gen_big_cnt_ic_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_big_cnt_ic_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_big_cnt_ic_cend <= io_job_job_0_big_cnt_ic_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_big_a <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_big_a <= io_job_job_0_big_a; // @[gen_addr.scala 293:11]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_max_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_max_addr <= io_job_job_0_small_0_max_addr; // @[gen_addr.scala 56:18]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_now_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_now_addr <= io_job_job_0_small_0_begin_addr; // @[gen_addr.scala 58:18]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (~state) begin // @[gen_addr.scala 266:18]
        gen_0_small_0_now_addr <= gen_small_0_y_begin_addr_nxt; // @[gen_addr.scala 266:18]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_cnt_ic_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (~state) begin // @[utils.scala 18:14]
        gen_0_small_0_cnt_ic_ccnt <= _gen_small_0_cnt_ic_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_cnt_ic_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_cnt_ic_cend <= io_job_job_0_small_0_cnt_ic_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_cnt_y_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_cnt_y_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_0_small_0_cnt_y_ccnt <= _GEN_38;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_cnt_y_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_cnt_y_cend <= io_job_job_0_small_0_cnt_y_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_bank_id <= 3'h0; // @[gen_addr.scala 64:17]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_0_small_0_bank_id <= _GEN_71;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_a <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_a <= io_job_job_0_small_0_a; // @[gen_addr.scala 271:11]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_ano_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_ano_bank_id <= io_job_job_0_small_0_ano_bank_id; // @[gen_addr.scala 272:21]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_0_small_0_ano_bank_id <= _GEN_73;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_cnt_swap_ccnt <= 1'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_cnt_swap_ccnt <= 1'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_0_small_0_cnt_swap_ccnt <= _GEN_66;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_cnt_swap_cend <= 1'h0; // @[write.scala 71:22]
    end else begin
      gen_0_small_0_cnt_swap_cend <= _GEN_214;
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_0_y_begin_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_0_y_begin_addr <= io_job_job_0_small_0_begin_addr; // @[gen_addr.scala 273:22]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_0_small_0_y_begin_addr <= _GEN_69;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_max_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_max_addr <= io_job_job_0_small_1_max_addr; // @[gen_addr.scala 56:18]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_now_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_now_addr <= io_job_job_0_small_1_begin_addr; // @[gen_addr.scala 58:18]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (~state) begin // @[gen_addr.scala 266:18]
        gen_0_small_1_now_addr <= gen_small_1_y_begin_addr_nxt; // @[gen_addr.scala 266:18]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_cnt_ic_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (~state) begin // @[utils.scala 18:14]
        gen_0_small_1_cnt_ic_ccnt <= _gen_small_1_cnt_ic_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_cnt_ic_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_cnt_ic_cend <= io_job_job_0_small_1_cnt_ic_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_cnt_y_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_cnt_y_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_0_small_1_cnt_y_ccnt <= _GEN_99;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_cnt_y_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_cnt_y_cend <= io_job_job_0_small_1_cnt_y_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_bank_id <= io_job_job_0_small_1_bank_id; // @[gen_addr.scala 64:17]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_0_small_1_bank_id <= _GEN_132;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_a <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_a <= io_job_job_0_small_1_a; // @[gen_addr.scala 271:11]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_ano_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_ano_bank_id <= io_job_job_0_small_1_ano_bank_id; // @[gen_addr.scala 272:21]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_0_small_1_ano_bank_id <= _GEN_134;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_cnt_swap_ccnt <= 1'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_cnt_swap_ccnt <= 1'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_0_small_1_cnt_swap_ccnt <= _GEN_127;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_cnt_swap_cend <= 1'h0; // @[write.scala 71:22]
    end else begin
      gen_0_small_1_cnt_swap_cend <= _GEN_231;
    end
    if (reset) begin // @[write.scala 71:22]
      gen_0_small_1_y_begin_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_0_small_1_y_begin_addr <= io_job_job_0_small_1_begin_addr; // @[gen_addr.scala 273:22]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_0_small_1_y_begin_addr <= _GEN_130;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_big_max_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_big_max_addr <= io_job_job_1_big_max_addr; // @[gen_addr.scala 56:18]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_big_now_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_big_now_addr <= io_job_job_1_big_begin_addr; // @[gen_addr.scala 58:18]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (state) begin // @[gen_addr.scala 288:18]
        gen_1_big_now_addr <= gen_big_now_addr_nxt; // @[gen_addr.scala 288:18]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_big_cnt_ic_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_big_cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (state) begin // @[utils.scala 18:14]
        gen_1_big_cnt_ic_ccnt <= _gen_big_cnt_ic_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_big_cnt_ic_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_big_cnt_ic_cend <= io_job_job_1_big_cnt_ic_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_big_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_big_bank_id <= io_job_job_1_big_bank_id; // @[gen_addr.scala 64:17]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_big_a <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_big_a <= io_job_job_1_big_a; // @[gen_addr.scala 293:11]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_max_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_max_addr <= io_job_job_1_small_0_max_addr; // @[gen_addr.scala 56:18]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_now_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_now_addr <= io_job_job_1_small_0_begin_addr; // @[gen_addr.scala 58:18]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (state) begin // @[gen_addr.scala 266:18]
        gen_1_small_0_now_addr <= gen_small_0_y_begin_addr_nxt; // @[gen_addr.scala 266:18]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_cnt_ic_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (state) begin // @[utils.scala 18:14]
        gen_1_small_0_cnt_ic_ccnt <= _gen_small_0_cnt_ic_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_cnt_ic_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_cnt_ic_cend <= io_job_job_1_small_0_cnt_ic_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_cnt_y_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_cnt_y_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_1_small_0_cnt_y_ccnt <= _GEN_39;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_cnt_y_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_cnt_y_cend <= io_job_job_1_small_0_cnt_y_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_bank_id <= io_job_job_1_small_0_bank_id; // @[gen_addr.scala 64:17]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_1_small_0_bank_id <= _GEN_72;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_a <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_a <= io_job_job_1_small_0_a; // @[gen_addr.scala 271:11]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_ano_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_ano_bank_id <= io_job_job_1_small_0_ano_bank_id; // @[gen_addr.scala 272:21]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_1_small_0_ano_bank_id <= _GEN_74;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_cnt_swap_ccnt <= 1'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_cnt_swap_ccnt <= 1'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_1_small_0_cnt_swap_ccnt <= _GEN_67;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_cnt_swap_cend <= 1'h0; // @[write.scala 71:22]
    end else begin
      gen_1_small_0_cnt_swap_cend <= _GEN_261;
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_0_y_begin_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_0_y_begin_addr <= io_job_job_1_small_0_begin_addr; // @[gen_addr.scala 273:22]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_1) begin // @[gen_addr.scala 250:27]
        gen_1_small_0_y_begin_addr <= _GEN_70;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_max_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_max_addr <= io_job_job_1_small_1_max_addr; // @[gen_addr.scala 56:18]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_now_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_now_addr <= io_job_job_1_small_1_begin_addr; // @[gen_addr.scala 58:18]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (state) begin // @[gen_addr.scala 266:18]
        gen_1_small_1_now_addr <= gen_small_1_y_begin_addr_nxt; // @[gen_addr.scala 266:18]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_cnt_ic_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (state) begin // @[utils.scala 18:14]
        gen_1_small_1_cnt_ic_ccnt <= _gen_small_1_cnt_ic_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_cnt_ic_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_cnt_ic_cend <= io_job_job_1_small_1_cnt_ic_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_cnt_y_ccnt <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_cnt_y_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_1_small_1_cnt_y_ccnt <= _GEN_100;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_cnt_y_cend <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_cnt_y_cend <= io_job_job_1_small_1_cnt_y_end; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_bank_id <= io_job_job_1_small_1_bank_id; // @[gen_addr.scala 64:17]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_1_small_1_bank_id <= _GEN_133;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_a <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_a <= io_job_job_1_small_1_a; // @[gen_addr.scala 271:11]
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_ano_bank_id <= 3'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_ano_bank_id <= io_job_job_1_small_1_ano_bank_id; // @[gen_addr.scala 272:21]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_1_small_1_ano_bank_id <= _GEN_135;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_cnt_swap_ccnt <= 1'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_cnt_swap_ccnt <= 1'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_1_small_1_cnt_swap_ccnt <= _GEN_128;
      end
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_cnt_swap_cend <= 1'h0; // @[write.scala 71:22]
    end else begin
      gen_1_small_1_cnt_swap_cend <= _GEN_278;
    end
    if (reset) begin // @[write.scala 71:22]
      gen_1_small_1_y_begin_addr <= 10'h0; // @[write.scala 71:22]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      gen_1_small_1_y_begin_addr <= io_job_job_1_small_1_begin_addr; // @[gen_addr.scala 273:22]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_4) begin // @[gen_addr.scala 250:27]
        gen_1_small_1_y_begin_addr <= _GEN_131;
      end
    end
    if (reset) begin // @[write.scala 72:25]
      cnt_ic_ccnt <= 10'h0; // @[write.scala 72:25]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      cnt_ic_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (io_valid_in) begin // @[write.scala 90:26]
      if (nxt_7) begin // @[utils.scala 18:20]
        cnt_ic_ccnt <= 10'h0;
      end else begin
        cnt_ic_ccnt <= _cnt_ic_ccnt_T_1;
      end
    end
    if (reset) begin // @[write.scala 72:25]
      cnt_ic_cend <= 10'h0; // @[write.scala 72:25]
    end else if (io_flag_job) begin // @[write.scala 85:22]
      cnt_ic_cend <= io_job_out_chan; // @[utils.scala 22:14]
    end
    if (reset) begin // @[write.scala 73:24]
      state <= 1'h0; // @[write.scala 73:24]
    end else if (!(io_flag_job)) begin // @[write.scala 85:22]
      if (io_valid_in) begin // @[write.scala 90:26]
        if (nxt_7) begin // @[write.scala 93:31]
          state <= ~state; // @[write.scala 94:23]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  gen_0_big_max_addr = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  gen_0_big_now_addr = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  gen_0_big_cnt_ic_ccnt = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  gen_0_big_cnt_ic_cend = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  gen_0_big_a = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  gen_0_small_0_max_addr = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  gen_0_small_0_now_addr = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  gen_0_small_0_cnt_ic_ccnt = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  gen_0_small_0_cnt_ic_cend = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  gen_0_small_0_cnt_y_ccnt = _RAND_9[9:0];
  _RAND_10 = {1{`RANDOM}};
  gen_0_small_0_cnt_y_cend = _RAND_10[9:0];
  _RAND_11 = {1{`RANDOM}};
  gen_0_small_0_bank_id = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  gen_0_small_0_a = _RAND_12[9:0];
  _RAND_13 = {1{`RANDOM}};
  gen_0_small_0_ano_bank_id = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  gen_0_small_0_cnt_swap_ccnt = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  gen_0_small_0_cnt_swap_cend = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  gen_0_small_0_y_begin_addr = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  gen_0_small_1_max_addr = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  gen_0_small_1_now_addr = _RAND_18[9:0];
  _RAND_19 = {1{`RANDOM}};
  gen_0_small_1_cnt_ic_ccnt = _RAND_19[9:0];
  _RAND_20 = {1{`RANDOM}};
  gen_0_small_1_cnt_ic_cend = _RAND_20[9:0];
  _RAND_21 = {1{`RANDOM}};
  gen_0_small_1_cnt_y_ccnt = _RAND_21[9:0];
  _RAND_22 = {1{`RANDOM}};
  gen_0_small_1_cnt_y_cend = _RAND_22[9:0];
  _RAND_23 = {1{`RANDOM}};
  gen_0_small_1_bank_id = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  gen_0_small_1_a = _RAND_24[9:0];
  _RAND_25 = {1{`RANDOM}};
  gen_0_small_1_ano_bank_id = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  gen_0_small_1_cnt_swap_ccnt = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  gen_0_small_1_cnt_swap_cend = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  gen_0_small_1_y_begin_addr = _RAND_28[9:0];
  _RAND_29 = {1{`RANDOM}};
  gen_1_big_max_addr = _RAND_29[9:0];
  _RAND_30 = {1{`RANDOM}};
  gen_1_big_now_addr = _RAND_30[9:0];
  _RAND_31 = {1{`RANDOM}};
  gen_1_big_cnt_ic_ccnt = _RAND_31[9:0];
  _RAND_32 = {1{`RANDOM}};
  gen_1_big_cnt_ic_cend = _RAND_32[9:0];
  _RAND_33 = {1{`RANDOM}};
  gen_1_big_bank_id = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  gen_1_big_a = _RAND_34[9:0];
  _RAND_35 = {1{`RANDOM}};
  gen_1_small_0_max_addr = _RAND_35[9:0];
  _RAND_36 = {1{`RANDOM}};
  gen_1_small_0_now_addr = _RAND_36[9:0];
  _RAND_37 = {1{`RANDOM}};
  gen_1_small_0_cnt_ic_ccnt = _RAND_37[9:0];
  _RAND_38 = {1{`RANDOM}};
  gen_1_small_0_cnt_ic_cend = _RAND_38[9:0];
  _RAND_39 = {1{`RANDOM}};
  gen_1_small_0_cnt_y_ccnt = _RAND_39[9:0];
  _RAND_40 = {1{`RANDOM}};
  gen_1_small_0_cnt_y_cend = _RAND_40[9:0];
  _RAND_41 = {1{`RANDOM}};
  gen_1_small_0_bank_id = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  gen_1_small_0_a = _RAND_42[9:0];
  _RAND_43 = {1{`RANDOM}};
  gen_1_small_0_ano_bank_id = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  gen_1_small_0_cnt_swap_ccnt = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  gen_1_small_0_cnt_swap_cend = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  gen_1_small_0_y_begin_addr = _RAND_46[9:0];
  _RAND_47 = {1{`RANDOM}};
  gen_1_small_1_max_addr = _RAND_47[9:0];
  _RAND_48 = {1{`RANDOM}};
  gen_1_small_1_now_addr = _RAND_48[9:0];
  _RAND_49 = {1{`RANDOM}};
  gen_1_small_1_cnt_ic_ccnt = _RAND_49[9:0];
  _RAND_50 = {1{`RANDOM}};
  gen_1_small_1_cnt_ic_cend = _RAND_50[9:0];
  _RAND_51 = {1{`RANDOM}};
  gen_1_small_1_cnt_y_ccnt = _RAND_51[9:0];
  _RAND_52 = {1{`RANDOM}};
  gen_1_small_1_cnt_y_cend = _RAND_52[9:0];
  _RAND_53 = {1{`RANDOM}};
  gen_1_small_1_bank_id = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  gen_1_small_1_a = _RAND_54[9:0];
  _RAND_55 = {1{`RANDOM}};
  gen_1_small_1_ano_bank_id = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  gen_1_small_1_cnt_swap_ccnt = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  gen_1_small_1_cnt_swap_cend = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  gen_1_small_1_y_begin_addr = _RAND_58[9:0];
  _RAND_59 = {1{`RANDOM}};
  cnt_ic_ccnt = _RAND_59[9:0];
  _RAND_60 = {1{`RANDOM}};
  cnt_ic_cend = _RAND_60[9:0];
  _RAND_61 = {1{`RANDOM}};
  state = _RAND_61[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ROMWeight(
  input         clock,
  input  [13:0] io_addr,
  output [15:0] io_out_0,
  output [15:0] io_out_1,
  output [15:0] io_out_2,
  output [15:0] io_out_3,
  output [15:0] io_out_4,
  output [15:0] io_out_5,
  output [15:0] io_out_6,
  output [15:0] io_out_7,
  output [15:0] io_out_8
);
  wire [13:0] weight0_addra; // @[bram.scala 223:21]
  wire  weight0_clka; // @[bram.scala 223:21]
  wire [143:0] weight0_douta; // @[bram.scala 223:21]
  wire [143:0] _WIRE_1 = weight0_douta;
  weight0 weight0 ( // @[bram.scala 223:21]
    .addra(weight0_addra),
    .clka(weight0_clka),
    .douta(weight0_douta)
  );
  assign io_out_0 = _WIRE_1[15:0]; // @[bram.scala 226:33]
  assign io_out_1 = _WIRE_1[31:16]; // @[bram.scala 226:33]
  assign io_out_2 = _WIRE_1[47:32]; // @[bram.scala 226:33]
  assign io_out_3 = _WIRE_1[63:48]; // @[bram.scala 226:33]
  assign io_out_4 = _WIRE_1[79:64]; // @[bram.scala 226:33]
  assign io_out_5 = _WIRE_1[95:80]; // @[bram.scala 226:33]
  assign io_out_6 = _WIRE_1[111:96]; // @[bram.scala 226:33]
  assign io_out_7 = _WIRE_1[127:112]; // @[bram.scala 226:33]
  assign io_out_8 = _WIRE_1[143:128]; // @[bram.scala 226:33]
  assign weight0_addra = io_addr; // @[bram.scala 225:15]
  assign weight0_clka = clock; // @[bram.scala 224:14]
endmodule
module ROMBias(
  input         clock,
  input  [7:0]  io_addr,
  output [35:0] io_out
);
  wire [7:0] bias0_addra; // @[bram.scala 210:21]
  wire  bias0_clka; // @[bram.scala 210:21]
  wire [35:0] bias0_douta; // @[bram.scala 210:21]
  bias0 bias0 ( // @[bram.scala 210:21]
    .addra(bias0_addra),
    .clka(bias0_clka),
    .douta(bias0_douta)
  );
  assign io_out = bias0_douta; // @[bram.scala 213:25]
  assign bias0_addra = io_addr; // @[bram.scala 212:15]
  assign bias0_clka = clock; // @[bram.scala 211:14]
endmodule
module RAMGroup(
  input         clock,
  input         reset,
  input         io_rd_valid_in,
  output        io_rd_valid_out,
  input  [2:0]  io_rd_addr1_addrs_0_bank_id,
  input  [9:0]  io_rd_addr1_addrs_1_addr,
  input  [9:0]  io_rd_addr2_addrs_1_addr,
  output [15:0] io_rd_big_0_data_0,
  output [15:0] io_rd_big_0_data_1,
  output [15:0] io_rd_big_0_data_2,
  output [15:0] io_rd_big_0_data_3,
  output [15:0] io_rd_big_0_data_4,
  output [15:0] io_rd_big_0_data_5,
  output [15:0] io_rd_big_0_data_6,
  output [15:0] io_rd_big_0_data_7,
  output [15:0] io_rd_big_0_data_8,
  output [15:0] io_rd_big_0_data_9,
  output [15:0] io_rd_big_0_data_10,
  output [15:0] io_rd_big_0_data_11,
  output [15:0] io_rd_big_0_data_12,
  output [15:0] io_rd_big_0_data_13,
  output [15:0] io_rd_big_0_data_14,
  output [15:0] io_rd_big_0_data_15,
  output [15:0] io_rd_big_0_data_16,
  output [15:0] io_rd_big_0_data_17,
  output [15:0] io_rd_big_0_data_18,
  output [15:0] io_rd_big_0_data_19,
  output [15:0] io_rd_big_0_data_20,
  output [15:0] io_rd_big_0_data_21,
  output [15:0] io_rd_big_0_data_22,
  output [15:0] io_rd_big_0_data_23,
  output [15:0] io_rd_big_0_data_24,
  output [15:0] io_rd_big_0_data_25,
  output [15:0] io_rd_big_0_data_26,
  output [15:0] io_rd_big_0_data_27,
  output [15:0] io_rd_big_0_data_28,
  output [15:0] io_rd_big_0_data_29,
  output [15:0] io_rd_big_0_data_30,
  output [15:0] io_rd_big_0_data_31,
  output [15:0] io_rd_big_0_data_32,
  output [15:0] io_rd_big_0_data_33,
  output [15:0] io_rd_big_0_data_34,
  output [15:0] io_rd_big_0_data_35,
  output [15:0] io_rd_big_0_data_36,
  output [15:0] io_rd_big_0_data_37,
  output [15:0] io_rd_big_0_data_38,
  output [15:0] io_rd_big_0_data_39,
  output [15:0] io_rd_big_0_data_40,
  output [15:0] io_rd_big_0_data_41,
  output [15:0] io_rd_big_0_data_42,
  output [15:0] io_rd_big_0_data_43,
  output [15:0] io_rd_big_0_data_44,
  output [15:0] io_rd_big_0_data_45,
  output [15:0] io_rd_big_0_data_46,
  output [15:0] io_rd_big_0_data_47,
  output [15:0] io_rd_big_1_data_0,
  output [15:0] io_rd_big_1_data_1,
  output [15:0] io_rd_big_1_data_2,
  output [15:0] io_rd_big_1_data_3,
  output [15:0] io_rd_big_1_data_4,
  output [15:0] io_rd_big_1_data_5,
  output [15:0] io_rd_big_1_data_6,
  output [15:0] io_rd_big_1_data_7,
  output [15:0] io_rd_big_1_data_8,
  output [15:0] io_rd_big_1_data_9,
  output [15:0] io_rd_big_1_data_10,
  output [15:0] io_rd_big_1_data_11,
  output [15:0] io_rd_big_1_data_12,
  output [15:0] io_rd_big_1_data_13,
  output [15:0] io_rd_big_1_data_14,
  output [15:0] io_rd_big_1_data_15,
  output [15:0] io_rd_big_1_data_16,
  output [15:0] io_rd_big_1_data_17,
  output [15:0] io_rd_big_1_data_18,
  output [15:0] io_rd_big_1_data_19,
  output [15:0] io_rd_big_1_data_20,
  output [15:0] io_rd_big_1_data_21,
  output [15:0] io_rd_big_1_data_22,
  output [15:0] io_rd_big_1_data_23,
  output [15:0] io_rd_big_1_data_24,
  output [15:0] io_rd_big_1_data_25,
  output [15:0] io_rd_big_1_data_26,
  output [15:0] io_rd_big_1_data_27,
  output [15:0] io_rd_big_1_data_28,
  output [15:0] io_rd_big_1_data_29,
  output [15:0] io_rd_big_1_data_30,
  output [15:0] io_rd_big_1_data_31,
  output [15:0] io_rd_big_1_data_32,
  output [15:0] io_rd_big_1_data_33,
  output [15:0] io_rd_big_1_data_34,
  output [15:0] io_rd_big_1_data_35,
  output [15:0] io_rd_big_1_data_36,
  output [15:0] io_rd_big_1_data_37,
  output [15:0] io_rd_big_1_data_38,
  output [15:0] io_rd_big_1_data_39,
  output [15:0] io_rd_big_1_data_40,
  output [15:0] io_rd_big_1_data_41,
  output [15:0] io_rd_big_1_data_42,
  output [15:0] io_rd_big_1_data_43,
  output [15:0] io_rd_big_1_data_44,
  output [15:0] io_rd_big_1_data_45,
  output [15:0] io_rd_big_1_data_46,
  output [15:0] io_rd_big_1_data_47,
  output [15:0] io_rd_small_0_0_data_0,
  output [15:0] io_rd_small_0_0_data_1,
  output [15:0] io_rd_small_0_0_data_2,
  output [15:0] io_rd_small_0_0_data_3,
  output [15:0] io_rd_small_0_0_data_4,
  output [15:0] io_rd_small_0_0_data_5,
  output [15:0] io_rd_small_0_0_data_6,
  output [15:0] io_rd_small_0_0_data_7,
  output [15:0] io_rd_small_0_1_data_0,
  output [15:0] io_rd_small_0_1_data_1,
  output [15:0] io_rd_small_0_1_data_2,
  output [15:0] io_rd_small_0_1_data_3,
  output [15:0] io_rd_small_0_1_data_4,
  output [15:0] io_rd_small_0_1_data_5,
  output [15:0] io_rd_small_0_1_data_6,
  output [15:0] io_rd_small_0_1_data_7,
  output [15:0] io_rd_small_0_2_data_0,
  output [15:0] io_rd_small_0_2_data_1,
  output [15:0] io_rd_small_0_2_data_2,
  output [15:0] io_rd_small_0_2_data_3,
  output [15:0] io_rd_small_0_2_data_4,
  output [15:0] io_rd_small_0_2_data_5,
  output [15:0] io_rd_small_0_2_data_6,
  output [15:0] io_rd_small_0_2_data_7,
  output [15:0] io_rd_small_0_3_data_0,
  output [15:0] io_rd_small_0_3_data_1,
  output [15:0] io_rd_small_0_3_data_2,
  output [15:0] io_rd_small_0_3_data_3,
  output [15:0] io_rd_small_0_3_data_4,
  output [15:0] io_rd_small_0_3_data_5,
  output [15:0] io_rd_small_0_3_data_6,
  output [15:0] io_rd_small_0_3_data_7,
  output [15:0] io_rd_small_1_0_data_0,
  output [15:0] io_rd_small_1_0_data_1,
  output [15:0] io_rd_small_1_0_data_2,
  output [15:0] io_rd_small_1_0_data_3,
  output [15:0] io_rd_small_1_0_data_4,
  output [15:0] io_rd_small_1_0_data_5,
  output [15:0] io_rd_small_1_0_data_6,
  output [15:0] io_rd_small_1_0_data_7,
  output [15:0] io_rd_small_1_1_data_0,
  output [15:0] io_rd_small_1_1_data_1,
  output [15:0] io_rd_small_1_1_data_2,
  output [15:0] io_rd_small_1_1_data_3,
  output [15:0] io_rd_small_1_1_data_4,
  output [15:0] io_rd_small_1_1_data_5,
  output [15:0] io_rd_small_1_1_data_6,
  output [15:0] io_rd_small_1_1_data_7,
  output [15:0] io_rd_small_1_2_data_0,
  output [15:0] io_rd_small_1_2_data_1,
  output [15:0] io_rd_small_1_2_data_2,
  output [15:0] io_rd_small_1_2_data_3,
  output [15:0] io_rd_small_1_2_data_4,
  output [15:0] io_rd_small_1_2_data_5,
  output [15:0] io_rd_small_1_2_data_6,
  output [15:0] io_rd_small_1_2_data_7,
  output [15:0] io_rd_small_1_3_data_0,
  output [15:0] io_rd_small_1_3_data_1,
  output [15:0] io_rd_small_1_3_data_2,
  output [15:0] io_rd_small_1_3_data_3,
  output [15:0] io_rd_small_1_3_data_4,
  output [15:0] io_rd_small_1_3_data_5,
  output [15:0] io_rd_small_1_3_data_6,
  output [15:0] io_rd_small_1_3_data_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [9:0] bram_big_bank0_addra; // @[bram.scala 96:27]
  wire  bram_big_bank0_clka; // @[bram.scala 96:27]
  wire [767:0] bram_big_bank0_dina; // @[bram.scala 96:27]
  wire [767:0] bram_big_bank0_douta; // @[bram.scala 96:27]
  wire  bram_big_bank0_wea; // @[bram.scala 96:27]
  wire [9:0] bram_big_bank0_addrb; // @[bram.scala 96:27]
  wire  bram_big_bank0_clkb; // @[bram.scala 96:27]
  wire [767:0] bram_big_bank0_dinb; // @[bram.scala 96:27]
  wire [767:0] bram_big_bank0_doutb; // @[bram.scala 96:27]
  wire  bram_big_bank0_web; // @[bram.scala 96:27]
  wire [9:0] bram_big_bank0_1_addra; // @[bram.scala 97:27]
  wire  bram_big_bank0_1_clka; // @[bram.scala 97:27]
  wire [767:0] bram_big_bank0_1_dina; // @[bram.scala 97:27]
  wire [767:0] bram_big_bank0_1_douta; // @[bram.scala 97:27]
  wire  bram_big_bank0_1_wea; // @[bram.scala 97:27]
  wire [9:0] bram_big_bank0_1_addrb; // @[bram.scala 97:27]
  wire  bram_big_bank0_1_clkb; // @[bram.scala 97:27]
  wire [767:0] bram_big_bank0_1_dinb; // @[bram.scala 97:27]
  wire [767:0] bram_big_bank0_1_doutb; // @[bram.scala 97:27]
  wire  bram_big_bank0_1_web; // @[bram.scala 97:27]
  wire [8:0] bram_small_bank0_addra; // @[bram.scala 99:29]
  wire  bram_small_bank0_clka; // @[bram.scala 99:29]
  wire [127:0] bram_small_bank0_dina; // @[bram.scala 99:29]
  wire [127:0] bram_small_bank0_douta; // @[bram.scala 99:29]
  wire  bram_small_bank0_wea; // @[bram.scala 99:29]
  wire [8:0] bram_small_bank0_addrb; // @[bram.scala 99:29]
  wire  bram_small_bank0_clkb; // @[bram.scala 99:29]
  wire [127:0] bram_small_bank0_dinb; // @[bram.scala 99:29]
  wire [127:0] bram_small_bank0_doutb; // @[bram.scala 99:29]
  wire  bram_small_bank0_web; // @[bram.scala 99:29]
  wire [8:0] bram_small_bank1_addra; // @[bram.scala 100:29]
  wire  bram_small_bank1_clka; // @[bram.scala 100:29]
  wire [127:0] bram_small_bank1_dina; // @[bram.scala 100:29]
  wire [127:0] bram_small_bank1_douta; // @[bram.scala 100:29]
  wire  bram_small_bank1_wea; // @[bram.scala 100:29]
  wire [8:0] bram_small_bank1_addrb; // @[bram.scala 100:29]
  wire  bram_small_bank1_clkb; // @[bram.scala 100:29]
  wire [127:0] bram_small_bank1_dinb; // @[bram.scala 100:29]
  wire [127:0] bram_small_bank1_doutb; // @[bram.scala 100:29]
  wire  bram_small_bank1_web; // @[bram.scala 100:29]
  wire [8:0] bram_small_bank2_addra; // @[bram.scala 101:29]
  wire  bram_small_bank2_clka; // @[bram.scala 101:29]
  wire [127:0] bram_small_bank2_dina; // @[bram.scala 101:29]
  wire [127:0] bram_small_bank2_douta; // @[bram.scala 101:29]
  wire  bram_small_bank2_wea; // @[bram.scala 101:29]
  wire [8:0] bram_small_bank2_addrb; // @[bram.scala 101:29]
  wire  bram_small_bank2_clkb; // @[bram.scala 101:29]
  wire [127:0] bram_small_bank2_dinb; // @[bram.scala 101:29]
  wire [127:0] bram_small_bank2_doutb; // @[bram.scala 101:29]
  wire  bram_small_bank2_web; // @[bram.scala 101:29]
  wire [8:0] bram_small_bank3_addra; // @[bram.scala 102:29]
  wire  bram_small_bank3_clka; // @[bram.scala 102:29]
  wire [127:0] bram_small_bank3_dina; // @[bram.scala 102:29]
  wire [127:0] bram_small_bank3_douta; // @[bram.scala 102:29]
  wire  bram_small_bank3_wea; // @[bram.scala 102:29]
  wire [8:0] bram_small_bank3_addrb; // @[bram.scala 102:29]
  wire  bram_small_bank3_clkb; // @[bram.scala 102:29]
  wire [127:0] bram_small_bank3_dinb; // @[bram.scala 102:29]
  wire [127:0] bram_small_bank3_doutb; // @[bram.scala 102:29]
  wire  bram_small_bank3_web; // @[bram.scala 102:29]
  wire [8:0] bram_small_bank4_addra; // @[bram.scala 103:29]
  wire  bram_small_bank4_clka; // @[bram.scala 103:29]
  wire [127:0] bram_small_bank4_dina; // @[bram.scala 103:29]
  wire [127:0] bram_small_bank4_douta; // @[bram.scala 103:29]
  wire  bram_small_bank4_wea; // @[bram.scala 103:29]
  wire [8:0] bram_small_bank4_addrb; // @[bram.scala 103:29]
  wire  bram_small_bank4_clkb; // @[bram.scala 103:29]
  wire [127:0] bram_small_bank4_dinb; // @[bram.scala 103:29]
  wire [127:0] bram_small_bank4_doutb; // @[bram.scala 103:29]
  wire  bram_small_bank4_web; // @[bram.scala 103:29]
  wire [8:0] bram_small_bank5_addra; // @[bram.scala 104:29]
  wire  bram_small_bank5_clka; // @[bram.scala 104:29]
  wire [127:0] bram_small_bank5_dina; // @[bram.scala 104:29]
  wire [127:0] bram_small_bank5_douta; // @[bram.scala 104:29]
  wire  bram_small_bank5_wea; // @[bram.scala 104:29]
  wire [8:0] bram_small_bank5_addrb; // @[bram.scala 104:29]
  wire  bram_small_bank5_clkb; // @[bram.scala 104:29]
  wire [127:0] bram_small_bank5_dinb; // @[bram.scala 104:29]
  wire [127:0] bram_small_bank5_doutb; // @[bram.scala 104:29]
  wire  bram_small_bank5_web; // @[bram.scala 104:29]
  wire [8:0] bram_small_bank6_addra; // @[bram.scala 105:29]
  wire  bram_small_bank6_clka; // @[bram.scala 105:29]
  wire [127:0] bram_small_bank6_dina; // @[bram.scala 105:29]
  wire [127:0] bram_small_bank6_douta; // @[bram.scala 105:29]
  wire  bram_small_bank6_wea; // @[bram.scala 105:29]
  wire [8:0] bram_small_bank6_addrb; // @[bram.scala 105:29]
  wire  bram_small_bank6_clkb; // @[bram.scala 105:29]
  wire [127:0] bram_small_bank6_dinb; // @[bram.scala 105:29]
  wire [127:0] bram_small_bank6_doutb; // @[bram.scala 105:29]
  wire  bram_small_bank6_web; // @[bram.scala 105:29]
  wire [8:0] bram_small_bank7_addra; // @[bram.scala 106:29]
  wire  bram_small_bank7_clka; // @[bram.scala 106:29]
  wire [127:0] bram_small_bank7_dina; // @[bram.scala 106:29]
  wire [127:0] bram_small_bank7_douta; // @[bram.scala 106:29]
  wire  bram_small_bank7_wea; // @[bram.scala 106:29]
  wire [8:0] bram_small_bank7_addrb; // @[bram.scala 106:29]
  wire  bram_small_bank7_clkb; // @[bram.scala 106:29]
  wire [127:0] bram_small_bank7_dinb; // @[bram.scala 106:29]
  wire [127:0] bram_small_bank7_doutb; // @[bram.scala 106:29]
  wire  bram_small_bank7_web; // @[bram.scala 106:29]
  reg  reg_valid; // @[bram.scala 87:28]
  reg  big_typ; // @[bram.scala 122:26]
  wire  _T_160 = io_rd_addr1_addrs_0_bank_id == 3'h0; // @[bram.scala 124:38]
  wire [767:0] big_banks_0_douta = bram_big_bank0_douta; // @[bram.scala 93:25 bram.scala 96:18]
  wire [15:0] _io_rd_big_0_T_1 = big_banks_0_douta[15:0]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_3 = big_banks_0_douta[31:16]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_5 = big_banks_0_douta[47:32]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_7 = big_banks_0_douta[63:48]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_9 = big_banks_0_douta[79:64]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_11 = big_banks_0_douta[95:80]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_13 = big_banks_0_douta[111:96]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_15 = big_banks_0_douta[127:112]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_17 = big_banks_0_douta[143:128]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_19 = big_banks_0_douta[159:144]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_21 = big_banks_0_douta[175:160]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_23 = big_banks_0_douta[191:176]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_25 = big_banks_0_douta[207:192]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_27 = big_banks_0_douta[223:208]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_29 = big_banks_0_douta[239:224]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_31 = big_banks_0_douta[255:240]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_33 = big_banks_0_douta[271:256]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_35 = big_banks_0_douta[287:272]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_37 = big_banks_0_douta[303:288]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_39 = big_banks_0_douta[319:304]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_41 = big_banks_0_douta[335:320]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_43 = big_banks_0_douta[351:336]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_45 = big_banks_0_douta[367:352]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_47 = big_banks_0_douta[383:368]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_49 = big_banks_0_douta[399:384]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_51 = big_banks_0_douta[415:400]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_53 = big_banks_0_douta[431:416]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_55 = big_banks_0_douta[447:432]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_57 = big_banks_0_douta[463:448]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_59 = big_banks_0_douta[479:464]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_61 = big_banks_0_douta[495:480]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_63 = big_banks_0_douta[511:496]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_65 = big_banks_0_douta[527:512]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_67 = big_banks_0_douta[543:528]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_69 = big_banks_0_douta[559:544]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_71 = big_banks_0_douta[575:560]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_73 = big_banks_0_douta[591:576]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_75 = big_banks_0_douta[607:592]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_77 = big_banks_0_douta[623:608]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_79 = big_banks_0_douta[639:624]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_81 = big_banks_0_douta[655:640]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_83 = big_banks_0_douta[671:656]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_85 = big_banks_0_douta[687:672]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_87 = big_banks_0_douta[703:688]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_89 = big_banks_0_douta[719:704]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_91 = big_banks_0_douta[735:720]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_93 = big_banks_0_douta[751:736]; // @[bram.scala 135:52]
  wire [15:0] _io_rd_big_0_T_95 = big_banks_0_douta[767:752]; // @[bram.scala 135:52]
  wire [767:0] big_banks_1_douta = bram_big_bank0_1_douta; // @[bram.scala 93:25 bram.scala 97:18]
  wire [15:0] _io_rd_big_1_T_1 = big_banks_1_douta[15:0]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_3 = big_banks_1_douta[31:16]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_5 = big_banks_1_douta[47:32]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_7 = big_banks_1_douta[63:48]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_9 = big_banks_1_douta[79:64]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_11 = big_banks_1_douta[95:80]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_13 = big_banks_1_douta[111:96]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_15 = big_banks_1_douta[127:112]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_17 = big_banks_1_douta[143:128]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_19 = big_banks_1_douta[159:144]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_21 = big_banks_1_douta[175:160]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_23 = big_banks_1_douta[191:176]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_25 = big_banks_1_douta[207:192]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_27 = big_banks_1_douta[223:208]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_29 = big_banks_1_douta[239:224]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_31 = big_banks_1_douta[255:240]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_33 = big_banks_1_douta[271:256]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_35 = big_banks_1_douta[287:272]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_37 = big_banks_1_douta[303:288]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_39 = big_banks_1_douta[319:304]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_41 = big_banks_1_douta[335:320]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_43 = big_banks_1_douta[351:336]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_45 = big_banks_1_douta[367:352]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_47 = big_banks_1_douta[383:368]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_49 = big_banks_1_douta[399:384]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_51 = big_banks_1_douta[415:400]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_53 = big_banks_1_douta[431:416]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_55 = big_banks_1_douta[447:432]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_57 = big_banks_1_douta[463:448]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_59 = big_banks_1_douta[479:464]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_61 = big_banks_1_douta[495:480]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_63 = big_banks_1_douta[511:496]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_65 = big_banks_1_douta[527:512]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_67 = big_banks_1_douta[543:528]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_69 = big_banks_1_douta[559:544]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_71 = big_banks_1_douta[575:560]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_73 = big_banks_1_douta[591:576]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_75 = big_banks_1_douta[607:592]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_77 = big_banks_1_douta[623:608]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_79 = big_banks_1_douta[639:624]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_81 = big_banks_1_douta[655:640]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_83 = big_banks_1_douta[671:656]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_85 = big_banks_1_douta[687:672]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_87 = big_banks_1_douta[703:688]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_89 = big_banks_1_douta[719:704]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_91 = big_banks_1_douta[735:720]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_93 = big_banks_1_douta[751:736]; // @[bram.scala 136:52]
  wire [15:0] _io_rd_big_1_T_95 = big_banks_1_douta[767:752]; // @[bram.scala 136:52]
  reg [1:0] typ_0; // @[bram.scala 143:22]
  reg [1:0] typ_1; // @[bram.scala 143:22]
  wire  _io_rd_small_0_0_T_8 = typ_0 == 2'h0; // @[bram.scala 171:26]
  wire [127:0] small_banks_0_douta = bram_small_bank0_douta; // @[bram.scala 94:27 bram.scala 99:20]
  wire [15:0] _io_rd_small_0_0_T_10 = small_banks_0_douta[15:0]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_12 = small_banks_0_douta[31:16]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_14 = small_banks_0_douta[47:32]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_16 = small_banks_0_douta[63:48]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_18 = small_banks_0_douta[79:64]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_20 = small_banks_0_douta[95:80]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_22 = small_banks_0_douta[111:96]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_24 = small_banks_0_douta[127:112]; // @[bram.scala 171:84]
  wire  _io_rd_small_0_0_T_25 = typ_0 == 2'h1; // @[bram.scala 171:26]
  wire [127:0] small_banks_1_douta = bram_small_bank1_douta; // @[bram.scala 94:27 bram.scala 100:20]
  wire [15:0] _io_rd_small_0_0_T_27 = small_banks_1_douta[15:0]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_29 = small_banks_1_douta[31:16]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_31 = small_banks_1_douta[47:32]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_33 = small_banks_1_douta[63:48]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_35 = small_banks_1_douta[79:64]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_37 = small_banks_1_douta[95:80]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_39 = small_banks_1_douta[111:96]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_41 = small_banks_1_douta[127:112]; // @[bram.scala 171:84]
  wire  _io_rd_small_0_0_T_42 = typ_0 == 2'h2; // @[bram.scala 171:26]
  wire [127:0] small_banks_2_douta = bram_small_bank2_douta; // @[bram.scala 94:27 bram.scala 101:20]
  wire [15:0] _io_rd_small_0_0_T_44 = small_banks_2_douta[15:0]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_46 = small_banks_2_douta[31:16]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_48 = small_banks_2_douta[47:32]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_50 = small_banks_2_douta[63:48]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_52 = small_banks_2_douta[79:64]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_54 = small_banks_2_douta[95:80]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_56 = small_banks_2_douta[111:96]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_58 = small_banks_2_douta[127:112]; // @[bram.scala 171:84]
  wire  _io_rd_small_0_0_T_59 = typ_0 == 2'h3; // @[bram.scala 171:26]
  wire [127:0] small_banks_3_douta = bram_small_bank3_douta; // @[bram.scala 94:27 bram.scala 102:20]
  wire [15:0] _io_rd_small_0_0_T_61 = small_banks_3_douta[15:0]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_63 = small_banks_3_douta[31:16]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_65 = small_banks_3_douta[47:32]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_67 = small_banks_3_douta[63:48]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_69 = small_banks_3_douta[79:64]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_71 = small_banks_3_douta[95:80]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_73 = small_banks_3_douta[111:96]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_75 = small_banks_3_douta[127:112]; // @[bram.scala 171:84]
  wire [15:0] _io_rd_small_0_0_T_76_data_0 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_61) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_76_data_1 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_63) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_76_data_2 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_65) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_76_data_3 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_67) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_76_data_4 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_69) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_76_data_5 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_71) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_76_data_6 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_73) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_76_data_7 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_75) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_77_data_0 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_44) : $signed(
    _io_rd_small_0_0_T_76_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_77_data_1 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_46) : $signed(
    _io_rd_small_0_0_T_76_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_77_data_2 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_48) : $signed(
    _io_rd_small_0_0_T_76_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_77_data_3 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_50) : $signed(
    _io_rd_small_0_0_T_76_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_77_data_4 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_52) : $signed(
    _io_rd_small_0_0_T_76_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_77_data_5 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_54) : $signed(
    _io_rd_small_0_0_T_76_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_77_data_6 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_56) : $signed(
    _io_rd_small_0_0_T_76_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_77_data_7 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_58) : $signed(
    _io_rd_small_0_0_T_76_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_78_data_0 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_27) : $signed(
    _io_rd_small_0_0_T_77_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_78_data_1 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_29) : $signed(
    _io_rd_small_0_0_T_77_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_78_data_2 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_31) : $signed(
    _io_rd_small_0_0_T_77_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_78_data_3 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_33) : $signed(
    _io_rd_small_0_0_T_77_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_78_data_4 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_35) : $signed(
    _io_rd_small_0_0_T_77_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_78_data_5 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_37) : $signed(
    _io_rd_small_0_0_T_77_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_78_data_6 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_39) : $signed(
    _io_rd_small_0_0_T_77_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_0_T_78_data_7 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_41) : $signed(
    _io_rd_small_0_0_T_77_data_7); // @[Mux.scala 98:16]
  wire [2:0] _GEN_125 = {{1'd0}, typ_1}; // @[bram.scala 174:26]
  wire  _io_rd_small_1_0_T_8 = _GEN_125 == 3'h4; // @[bram.scala 174:26]
  wire [127:0] small_banks_4_douta = bram_small_bank4_douta; // @[bram.scala 94:27 bram.scala 103:20]
  wire [15:0] _io_rd_small_1_0_T_10 = small_banks_4_douta[15:0]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_12 = small_banks_4_douta[31:16]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_14 = small_banks_4_douta[47:32]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_16 = small_banks_4_douta[63:48]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_18 = small_banks_4_douta[79:64]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_20 = small_banks_4_douta[95:80]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_22 = small_banks_4_douta[111:96]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_24 = small_banks_4_douta[127:112]; // @[bram.scala 174:90]
  wire  _io_rd_small_1_0_T_25 = _GEN_125 == 3'h5; // @[bram.scala 174:26]
  wire [127:0] small_banks_5_douta = bram_small_bank5_douta; // @[bram.scala 94:27 bram.scala 104:20]
  wire [15:0] _io_rd_small_1_0_T_27 = small_banks_5_douta[15:0]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_29 = small_banks_5_douta[31:16]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_31 = small_banks_5_douta[47:32]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_33 = small_banks_5_douta[63:48]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_35 = small_banks_5_douta[79:64]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_37 = small_banks_5_douta[95:80]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_39 = small_banks_5_douta[111:96]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_41 = small_banks_5_douta[127:112]; // @[bram.scala 174:90]
  wire  _io_rd_small_1_0_T_42 = _GEN_125 == 3'h6; // @[bram.scala 174:26]
  wire [127:0] small_banks_6_douta = bram_small_bank6_douta; // @[bram.scala 94:27 bram.scala 105:20]
  wire [15:0] _io_rd_small_1_0_T_44 = small_banks_6_douta[15:0]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_46 = small_banks_6_douta[31:16]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_48 = small_banks_6_douta[47:32]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_50 = small_banks_6_douta[63:48]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_52 = small_banks_6_douta[79:64]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_54 = small_banks_6_douta[95:80]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_56 = small_banks_6_douta[111:96]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_58 = small_banks_6_douta[127:112]; // @[bram.scala 174:90]
  wire  _io_rd_small_1_0_T_59 = _GEN_125 == 3'h7; // @[bram.scala 174:26]
  wire [127:0] small_banks_7_douta = bram_small_bank7_douta; // @[bram.scala 94:27 bram.scala 106:20]
  wire [15:0] _io_rd_small_1_0_T_61 = small_banks_7_douta[15:0]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_63 = small_banks_7_douta[31:16]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_65 = small_banks_7_douta[47:32]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_67 = small_banks_7_douta[63:48]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_69 = small_banks_7_douta[79:64]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_71 = small_banks_7_douta[95:80]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_73 = small_banks_7_douta[111:96]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_75 = small_banks_7_douta[127:112]; // @[bram.scala 174:90]
  wire [15:0] _io_rd_small_1_0_T_76_data_0 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_61) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_76_data_1 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_63) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_76_data_2 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_65) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_76_data_3 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_67) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_76_data_4 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_69) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_76_data_5 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_71) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_76_data_6 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_73) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_76_data_7 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_75) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_77_data_0 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_44) : $signed(
    _io_rd_small_1_0_T_76_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_77_data_1 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_46) : $signed(
    _io_rd_small_1_0_T_76_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_77_data_2 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_48) : $signed(
    _io_rd_small_1_0_T_76_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_77_data_3 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_50) : $signed(
    _io_rd_small_1_0_T_76_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_77_data_4 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_52) : $signed(
    _io_rd_small_1_0_T_76_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_77_data_5 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_54) : $signed(
    _io_rd_small_1_0_T_76_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_77_data_6 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_56) : $signed(
    _io_rd_small_1_0_T_76_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_77_data_7 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_58) : $signed(
    _io_rd_small_1_0_T_76_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_78_data_0 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_27) : $signed(
    _io_rd_small_1_0_T_77_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_78_data_1 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_29) : $signed(
    _io_rd_small_1_0_T_77_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_78_data_2 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_31) : $signed(
    _io_rd_small_1_0_T_77_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_78_data_3 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_33) : $signed(
    _io_rd_small_1_0_T_77_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_78_data_4 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_35) : $signed(
    _io_rd_small_1_0_T_77_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_78_data_5 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_37) : $signed(
    _io_rd_small_1_0_T_77_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_78_data_6 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_39) : $signed(
    _io_rd_small_1_0_T_77_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_0_T_78_data_7 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_41) : $signed(
    _io_rd_small_1_0_T_77_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_76_data_0 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_10) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_76_data_1 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_12) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_76_data_2 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_14) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_76_data_3 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_16) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_76_data_4 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_18) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_76_data_5 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_20) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_76_data_6 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_22) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_76_data_7 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_24) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_77_data_0 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_61) : $signed(
    _io_rd_small_0_1_T_76_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_77_data_1 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_63) : $signed(
    _io_rd_small_0_1_T_76_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_77_data_2 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_65) : $signed(
    _io_rd_small_0_1_T_76_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_77_data_3 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_67) : $signed(
    _io_rd_small_0_1_T_76_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_77_data_4 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_69) : $signed(
    _io_rd_small_0_1_T_76_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_77_data_5 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_71) : $signed(
    _io_rd_small_0_1_T_76_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_77_data_6 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_73) : $signed(
    _io_rd_small_0_1_T_76_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_77_data_7 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_75) : $signed(
    _io_rd_small_0_1_T_76_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_78_data_0 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_44) : $signed(
    _io_rd_small_0_1_T_77_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_78_data_1 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_46) : $signed(
    _io_rd_small_0_1_T_77_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_78_data_2 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_48) : $signed(
    _io_rd_small_0_1_T_77_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_78_data_3 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_50) : $signed(
    _io_rd_small_0_1_T_77_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_78_data_4 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_52) : $signed(
    _io_rd_small_0_1_T_77_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_78_data_5 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_54) : $signed(
    _io_rd_small_0_1_T_77_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_78_data_6 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_56) : $signed(
    _io_rd_small_0_1_T_77_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_1_T_78_data_7 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_58) : $signed(
    _io_rd_small_0_1_T_77_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_76_data_0 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_10) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_76_data_1 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_12) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_76_data_2 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_14) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_76_data_3 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_16) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_76_data_4 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_18) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_76_data_5 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_20) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_76_data_6 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_22) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_76_data_7 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_24) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_77_data_0 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_61) : $signed(
    _io_rd_small_1_1_T_76_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_77_data_1 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_63) : $signed(
    _io_rd_small_1_1_T_76_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_77_data_2 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_65) : $signed(
    _io_rd_small_1_1_T_76_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_77_data_3 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_67) : $signed(
    _io_rd_small_1_1_T_76_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_77_data_4 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_69) : $signed(
    _io_rd_small_1_1_T_76_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_77_data_5 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_71) : $signed(
    _io_rd_small_1_1_T_76_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_77_data_6 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_73) : $signed(
    _io_rd_small_1_1_T_76_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_77_data_7 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_75) : $signed(
    _io_rd_small_1_1_T_76_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_78_data_0 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_44) : $signed(
    _io_rd_small_1_1_T_77_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_78_data_1 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_46) : $signed(
    _io_rd_small_1_1_T_77_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_78_data_2 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_48) : $signed(
    _io_rd_small_1_1_T_77_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_78_data_3 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_50) : $signed(
    _io_rd_small_1_1_T_77_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_78_data_4 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_52) : $signed(
    _io_rd_small_1_1_T_77_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_78_data_5 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_54) : $signed(
    _io_rd_small_1_1_T_77_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_78_data_6 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_56) : $signed(
    _io_rd_small_1_1_T_77_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_1_T_78_data_7 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_58) : $signed(
    _io_rd_small_1_1_T_77_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_76_data_0 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_27) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_76_data_1 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_29) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_76_data_2 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_31) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_76_data_3 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_33) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_76_data_4 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_35) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_76_data_5 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_37) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_76_data_6 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_39) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_76_data_7 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_41) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_77_data_0 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_10) : $signed(
    _io_rd_small_0_2_T_76_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_77_data_1 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_12) : $signed(
    _io_rd_small_0_2_T_76_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_77_data_2 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_14) : $signed(
    _io_rd_small_0_2_T_76_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_77_data_3 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_16) : $signed(
    _io_rd_small_0_2_T_76_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_77_data_4 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_18) : $signed(
    _io_rd_small_0_2_T_76_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_77_data_5 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_20) : $signed(
    _io_rd_small_0_2_T_76_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_77_data_6 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_22) : $signed(
    _io_rd_small_0_2_T_76_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_77_data_7 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_24) : $signed(
    _io_rd_small_0_2_T_76_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_78_data_0 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_61) : $signed(
    _io_rd_small_0_2_T_77_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_78_data_1 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_63) : $signed(
    _io_rd_small_0_2_T_77_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_78_data_2 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_65) : $signed(
    _io_rd_small_0_2_T_77_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_78_data_3 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_67) : $signed(
    _io_rd_small_0_2_T_77_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_78_data_4 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_69) : $signed(
    _io_rd_small_0_2_T_77_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_78_data_5 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_71) : $signed(
    _io_rd_small_0_2_T_77_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_78_data_6 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_73) : $signed(
    _io_rd_small_0_2_T_77_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_2_T_78_data_7 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_75) : $signed(
    _io_rd_small_0_2_T_77_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_76_data_0 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_27) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_76_data_1 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_29) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_76_data_2 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_31) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_76_data_3 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_33) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_76_data_4 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_35) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_76_data_5 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_37) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_76_data_6 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_39) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_76_data_7 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_41) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_77_data_0 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_10) : $signed(
    _io_rd_small_1_2_T_76_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_77_data_1 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_12) : $signed(
    _io_rd_small_1_2_T_76_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_77_data_2 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_14) : $signed(
    _io_rd_small_1_2_T_76_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_77_data_3 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_16) : $signed(
    _io_rd_small_1_2_T_76_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_77_data_4 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_18) : $signed(
    _io_rd_small_1_2_T_76_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_77_data_5 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_20) : $signed(
    _io_rd_small_1_2_T_76_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_77_data_6 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_22) : $signed(
    _io_rd_small_1_2_T_76_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_77_data_7 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_24) : $signed(
    _io_rd_small_1_2_T_76_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_78_data_0 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_61) : $signed(
    _io_rd_small_1_2_T_77_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_78_data_1 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_63) : $signed(
    _io_rd_small_1_2_T_77_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_78_data_2 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_65) : $signed(
    _io_rd_small_1_2_T_77_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_78_data_3 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_67) : $signed(
    _io_rd_small_1_2_T_77_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_78_data_4 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_69) : $signed(
    _io_rd_small_1_2_T_77_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_78_data_5 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_71) : $signed(
    _io_rd_small_1_2_T_77_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_78_data_6 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_73) : $signed(
    _io_rd_small_1_2_T_77_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_2_T_78_data_7 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_75) : $signed(
    _io_rd_small_1_2_T_77_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_76_data_0 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_44) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_76_data_1 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_46) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_76_data_2 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_48) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_76_data_3 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_50) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_76_data_4 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_52) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_76_data_5 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_54) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_76_data_6 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_56) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_76_data_7 = _io_rd_small_0_0_T_59 ? $signed(_io_rd_small_0_0_T_58) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_77_data_0 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_27) : $signed(
    _io_rd_small_0_3_T_76_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_77_data_1 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_29) : $signed(
    _io_rd_small_0_3_T_76_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_77_data_2 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_31) : $signed(
    _io_rd_small_0_3_T_76_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_77_data_3 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_33) : $signed(
    _io_rd_small_0_3_T_76_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_77_data_4 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_35) : $signed(
    _io_rd_small_0_3_T_76_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_77_data_5 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_37) : $signed(
    _io_rd_small_0_3_T_76_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_77_data_6 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_39) : $signed(
    _io_rd_small_0_3_T_76_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_77_data_7 = _io_rd_small_0_0_T_42 ? $signed(_io_rd_small_0_0_T_41) : $signed(
    _io_rd_small_0_3_T_76_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_78_data_0 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_10) : $signed(
    _io_rd_small_0_3_T_77_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_78_data_1 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_12) : $signed(
    _io_rd_small_0_3_T_77_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_78_data_2 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_14) : $signed(
    _io_rd_small_0_3_T_77_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_78_data_3 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_16) : $signed(
    _io_rd_small_0_3_T_77_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_78_data_4 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_18) : $signed(
    _io_rd_small_0_3_T_77_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_78_data_5 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_20) : $signed(
    _io_rd_small_0_3_T_77_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_78_data_6 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_22) : $signed(
    _io_rd_small_0_3_T_77_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_0_3_T_78_data_7 = _io_rd_small_0_0_T_25 ? $signed(_io_rd_small_0_0_T_24) : $signed(
    _io_rd_small_0_3_T_77_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_76_data_0 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_44) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_76_data_1 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_46) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_76_data_2 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_48) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_76_data_3 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_50) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_76_data_4 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_52) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_76_data_5 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_54) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_76_data_6 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_56) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_76_data_7 = _io_rd_small_1_0_T_59 ? $signed(_io_rd_small_1_0_T_58) : $signed(16'sh0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_77_data_0 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_27) : $signed(
    _io_rd_small_1_3_T_76_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_77_data_1 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_29) : $signed(
    _io_rd_small_1_3_T_76_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_77_data_2 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_31) : $signed(
    _io_rd_small_1_3_T_76_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_77_data_3 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_33) : $signed(
    _io_rd_small_1_3_T_76_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_77_data_4 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_35) : $signed(
    _io_rd_small_1_3_T_76_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_77_data_5 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_37) : $signed(
    _io_rd_small_1_3_T_76_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_77_data_6 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_39) : $signed(
    _io_rd_small_1_3_T_76_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_77_data_7 = _io_rd_small_1_0_T_42 ? $signed(_io_rd_small_1_0_T_41) : $signed(
    _io_rd_small_1_3_T_76_data_7); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_78_data_0 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_10) : $signed(
    _io_rd_small_1_3_T_77_data_0); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_78_data_1 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_12) : $signed(
    _io_rd_small_1_3_T_77_data_1); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_78_data_2 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_14) : $signed(
    _io_rd_small_1_3_T_77_data_2); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_78_data_3 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_16) : $signed(
    _io_rd_small_1_3_T_77_data_3); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_78_data_4 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_18) : $signed(
    _io_rd_small_1_3_T_77_data_4); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_78_data_5 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_20) : $signed(
    _io_rd_small_1_3_T_77_data_5); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_78_data_6 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_22) : $signed(
    _io_rd_small_1_3_T_77_data_6); // @[Mux.scala 98:16]
  wire [15:0] _io_rd_small_1_3_T_78_data_7 = _io_rd_small_1_0_T_25 ? $signed(_io_rd_small_1_0_T_24) : $signed(
    _io_rd_small_1_3_T_77_data_7); // @[Mux.scala 98:16]
  bram_big_bank0 bram_big_bank0 ( // @[bram.scala 96:27]
    .addra(bram_big_bank0_addra),
    .clka(bram_big_bank0_clka),
    .dina(bram_big_bank0_dina),
    .douta(bram_big_bank0_douta),
    .wea(bram_big_bank0_wea),
    .addrb(bram_big_bank0_addrb),
    .clkb(bram_big_bank0_clkb),
    .dinb(bram_big_bank0_dinb),
    .doutb(bram_big_bank0_doutb),
    .web(bram_big_bank0_web)
  );
  bram_big_bank0 bram_big_bank0_1 ( // @[bram.scala 97:27]
    .addra(bram_big_bank0_1_addra),
    .clka(bram_big_bank0_1_clka),
    .dina(bram_big_bank0_1_dina),
    .douta(bram_big_bank0_1_douta),
    .wea(bram_big_bank0_1_wea),
    .addrb(bram_big_bank0_1_addrb),
    .clkb(bram_big_bank0_1_clkb),
    .dinb(bram_big_bank0_1_dinb),
    .doutb(bram_big_bank0_1_doutb),
    .web(bram_big_bank0_1_web)
  );
  bram_small_bank0 bram_small_bank0 ( // @[bram.scala 99:29]
    .addra(bram_small_bank0_addra),
    .clka(bram_small_bank0_clka),
    .dina(bram_small_bank0_dina),
    .douta(bram_small_bank0_douta),
    .wea(bram_small_bank0_wea),
    .addrb(bram_small_bank0_addrb),
    .clkb(bram_small_bank0_clkb),
    .dinb(bram_small_bank0_dinb),
    .doutb(bram_small_bank0_doutb),
    .web(bram_small_bank0_web)
  );
  bram_small_bank1 bram_small_bank1 ( // @[bram.scala 100:29]
    .addra(bram_small_bank1_addra),
    .clka(bram_small_bank1_clka),
    .dina(bram_small_bank1_dina),
    .douta(bram_small_bank1_douta),
    .wea(bram_small_bank1_wea),
    .addrb(bram_small_bank1_addrb),
    .clkb(bram_small_bank1_clkb),
    .dinb(bram_small_bank1_dinb),
    .doutb(bram_small_bank1_doutb),
    .web(bram_small_bank1_web)
  );
  bram_small_bank2 bram_small_bank2 ( // @[bram.scala 101:29]
    .addra(bram_small_bank2_addra),
    .clka(bram_small_bank2_clka),
    .dina(bram_small_bank2_dina),
    .douta(bram_small_bank2_douta),
    .wea(bram_small_bank2_wea),
    .addrb(bram_small_bank2_addrb),
    .clkb(bram_small_bank2_clkb),
    .dinb(bram_small_bank2_dinb),
    .doutb(bram_small_bank2_doutb),
    .web(bram_small_bank2_web)
  );
  bram_small_bank3 bram_small_bank3 ( // @[bram.scala 102:29]
    .addra(bram_small_bank3_addra),
    .clka(bram_small_bank3_clka),
    .dina(bram_small_bank3_dina),
    .douta(bram_small_bank3_douta),
    .wea(bram_small_bank3_wea),
    .addrb(bram_small_bank3_addrb),
    .clkb(bram_small_bank3_clkb),
    .dinb(bram_small_bank3_dinb),
    .doutb(bram_small_bank3_doutb),
    .web(bram_small_bank3_web)
  );
  bram_small_bank4 bram_small_bank4 ( // @[bram.scala 103:29]
    .addra(bram_small_bank4_addra),
    .clka(bram_small_bank4_clka),
    .dina(bram_small_bank4_dina),
    .douta(bram_small_bank4_douta),
    .wea(bram_small_bank4_wea),
    .addrb(bram_small_bank4_addrb),
    .clkb(bram_small_bank4_clkb),
    .dinb(bram_small_bank4_dinb),
    .doutb(bram_small_bank4_doutb),
    .web(bram_small_bank4_web)
  );
  bram_small_bank5 bram_small_bank5 ( // @[bram.scala 104:29]
    .addra(bram_small_bank5_addra),
    .clka(bram_small_bank5_clka),
    .dina(bram_small_bank5_dina),
    .douta(bram_small_bank5_douta),
    .wea(bram_small_bank5_wea),
    .addrb(bram_small_bank5_addrb),
    .clkb(bram_small_bank5_clkb),
    .dinb(bram_small_bank5_dinb),
    .doutb(bram_small_bank5_doutb),
    .web(bram_small_bank5_web)
  );
  bram_small_bank6 bram_small_bank6 ( // @[bram.scala 105:29]
    .addra(bram_small_bank6_addra),
    .clka(bram_small_bank6_clka),
    .dina(bram_small_bank6_dina),
    .douta(bram_small_bank6_douta),
    .wea(bram_small_bank6_wea),
    .addrb(bram_small_bank6_addrb),
    .clkb(bram_small_bank6_clkb),
    .dinb(bram_small_bank6_dinb),
    .doutb(bram_small_bank6_doutb),
    .web(bram_small_bank6_web)
  );
  bram_small_bank7 bram_small_bank7 ( // @[bram.scala 106:29]
    .addra(bram_small_bank7_addra),
    .clka(bram_small_bank7_clka),
    .dina(bram_small_bank7_dina),
    .douta(bram_small_bank7_douta),
    .wea(bram_small_bank7_wea),
    .addrb(bram_small_bank7_addrb),
    .clkb(bram_small_bank7_clkb),
    .dinb(bram_small_bank7_dinb),
    .doutb(bram_small_bank7_doutb),
    .web(bram_small_bank7_web)
  );
  assign io_rd_valid_out = reg_valid; // @[bram.scala 88:21]
  assign io_rd_big_0_data_0 = big_typ ? $signed(_io_rd_big_0_T_1) : $signed(_io_rd_big_1_T_1); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_1 = big_typ ? $signed(_io_rd_big_0_T_3) : $signed(_io_rd_big_1_T_3); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_2 = big_typ ? $signed(_io_rd_big_0_T_5) : $signed(_io_rd_big_1_T_5); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_3 = big_typ ? $signed(_io_rd_big_0_T_7) : $signed(_io_rd_big_1_T_7); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_4 = big_typ ? $signed(_io_rd_big_0_T_9) : $signed(_io_rd_big_1_T_9); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_5 = big_typ ? $signed(_io_rd_big_0_T_11) : $signed(_io_rd_big_1_T_11); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_6 = big_typ ? $signed(_io_rd_big_0_T_13) : $signed(_io_rd_big_1_T_13); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_7 = big_typ ? $signed(_io_rd_big_0_T_15) : $signed(_io_rd_big_1_T_15); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_8 = big_typ ? $signed(_io_rd_big_0_T_17) : $signed(_io_rd_big_1_T_17); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_9 = big_typ ? $signed(_io_rd_big_0_T_19) : $signed(_io_rd_big_1_T_19); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_10 = big_typ ? $signed(_io_rd_big_0_T_21) : $signed(_io_rd_big_1_T_21); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_11 = big_typ ? $signed(_io_rd_big_0_T_23) : $signed(_io_rd_big_1_T_23); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_12 = big_typ ? $signed(_io_rd_big_0_T_25) : $signed(_io_rd_big_1_T_25); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_13 = big_typ ? $signed(_io_rd_big_0_T_27) : $signed(_io_rd_big_1_T_27); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_14 = big_typ ? $signed(_io_rd_big_0_T_29) : $signed(_io_rd_big_1_T_29); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_15 = big_typ ? $signed(_io_rd_big_0_T_31) : $signed(_io_rd_big_1_T_31); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_16 = big_typ ? $signed(_io_rd_big_0_T_33) : $signed(_io_rd_big_1_T_33); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_17 = big_typ ? $signed(_io_rd_big_0_T_35) : $signed(_io_rd_big_1_T_35); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_18 = big_typ ? $signed(_io_rd_big_0_T_37) : $signed(_io_rd_big_1_T_37); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_19 = big_typ ? $signed(_io_rd_big_0_T_39) : $signed(_io_rd_big_1_T_39); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_20 = big_typ ? $signed(_io_rd_big_0_T_41) : $signed(_io_rd_big_1_T_41); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_21 = big_typ ? $signed(_io_rd_big_0_T_43) : $signed(_io_rd_big_1_T_43); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_22 = big_typ ? $signed(_io_rd_big_0_T_45) : $signed(_io_rd_big_1_T_45); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_23 = big_typ ? $signed(_io_rd_big_0_T_47) : $signed(_io_rd_big_1_T_47); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_24 = big_typ ? $signed(_io_rd_big_0_T_49) : $signed(_io_rd_big_1_T_49); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_25 = big_typ ? $signed(_io_rd_big_0_T_51) : $signed(_io_rd_big_1_T_51); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_26 = big_typ ? $signed(_io_rd_big_0_T_53) : $signed(_io_rd_big_1_T_53); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_27 = big_typ ? $signed(_io_rd_big_0_T_55) : $signed(_io_rd_big_1_T_55); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_28 = big_typ ? $signed(_io_rd_big_0_T_57) : $signed(_io_rd_big_1_T_57); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_29 = big_typ ? $signed(_io_rd_big_0_T_59) : $signed(_io_rd_big_1_T_59); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_30 = big_typ ? $signed(_io_rd_big_0_T_61) : $signed(_io_rd_big_1_T_61); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_31 = big_typ ? $signed(_io_rd_big_0_T_63) : $signed(_io_rd_big_1_T_63); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_32 = big_typ ? $signed(_io_rd_big_0_T_65) : $signed(_io_rd_big_1_T_65); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_33 = big_typ ? $signed(_io_rd_big_0_T_67) : $signed(_io_rd_big_1_T_67); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_34 = big_typ ? $signed(_io_rd_big_0_T_69) : $signed(_io_rd_big_1_T_69); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_35 = big_typ ? $signed(_io_rd_big_0_T_71) : $signed(_io_rd_big_1_T_71); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_36 = big_typ ? $signed(_io_rd_big_0_T_73) : $signed(_io_rd_big_1_T_73); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_37 = big_typ ? $signed(_io_rd_big_0_T_75) : $signed(_io_rd_big_1_T_75); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_38 = big_typ ? $signed(_io_rd_big_0_T_77) : $signed(_io_rd_big_1_T_77); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_39 = big_typ ? $signed(_io_rd_big_0_T_79) : $signed(_io_rd_big_1_T_79); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_40 = big_typ ? $signed(_io_rd_big_0_T_81) : $signed(_io_rd_big_1_T_81); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_41 = big_typ ? $signed(_io_rd_big_0_T_83) : $signed(_io_rd_big_1_T_83); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_42 = big_typ ? $signed(_io_rd_big_0_T_85) : $signed(_io_rd_big_1_T_85); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_43 = big_typ ? $signed(_io_rd_big_0_T_87) : $signed(_io_rd_big_1_T_87); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_44 = big_typ ? $signed(_io_rd_big_0_T_89) : $signed(_io_rd_big_1_T_89); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_45 = big_typ ? $signed(_io_rd_big_0_T_91) : $signed(_io_rd_big_1_T_91); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_46 = big_typ ? $signed(_io_rd_big_0_T_93) : $signed(_io_rd_big_1_T_93); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_0_data_47 = big_typ ? $signed(_io_rd_big_0_T_95) : $signed(_io_rd_big_1_T_95); // @[bram.scala 134:24 bram.scala 135:22 bram.scala 139:22]
  assign io_rd_big_1_data_0 = big_typ ? $signed(_io_rd_big_1_T_1) : $signed(_io_rd_big_0_T_1); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_1 = big_typ ? $signed(_io_rd_big_1_T_3) : $signed(_io_rd_big_0_T_3); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_2 = big_typ ? $signed(_io_rd_big_1_T_5) : $signed(_io_rd_big_0_T_5); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_3 = big_typ ? $signed(_io_rd_big_1_T_7) : $signed(_io_rd_big_0_T_7); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_4 = big_typ ? $signed(_io_rd_big_1_T_9) : $signed(_io_rd_big_0_T_9); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_5 = big_typ ? $signed(_io_rd_big_1_T_11) : $signed(_io_rd_big_0_T_11); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_6 = big_typ ? $signed(_io_rd_big_1_T_13) : $signed(_io_rd_big_0_T_13); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_7 = big_typ ? $signed(_io_rd_big_1_T_15) : $signed(_io_rd_big_0_T_15); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_8 = big_typ ? $signed(_io_rd_big_1_T_17) : $signed(_io_rd_big_0_T_17); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_9 = big_typ ? $signed(_io_rd_big_1_T_19) : $signed(_io_rd_big_0_T_19); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_10 = big_typ ? $signed(_io_rd_big_1_T_21) : $signed(_io_rd_big_0_T_21); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_11 = big_typ ? $signed(_io_rd_big_1_T_23) : $signed(_io_rd_big_0_T_23); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_12 = big_typ ? $signed(_io_rd_big_1_T_25) : $signed(_io_rd_big_0_T_25); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_13 = big_typ ? $signed(_io_rd_big_1_T_27) : $signed(_io_rd_big_0_T_27); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_14 = big_typ ? $signed(_io_rd_big_1_T_29) : $signed(_io_rd_big_0_T_29); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_15 = big_typ ? $signed(_io_rd_big_1_T_31) : $signed(_io_rd_big_0_T_31); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_16 = big_typ ? $signed(_io_rd_big_1_T_33) : $signed(_io_rd_big_0_T_33); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_17 = big_typ ? $signed(_io_rd_big_1_T_35) : $signed(_io_rd_big_0_T_35); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_18 = big_typ ? $signed(_io_rd_big_1_T_37) : $signed(_io_rd_big_0_T_37); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_19 = big_typ ? $signed(_io_rd_big_1_T_39) : $signed(_io_rd_big_0_T_39); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_20 = big_typ ? $signed(_io_rd_big_1_T_41) : $signed(_io_rd_big_0_T_41); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_21 = big_typ ? $signed(_io_rd_big_1_T_43) : $signed(_io_rd_big_0_T_43); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_22 = big_typ ? $signed(_io_rd_big_1_T_45) : $signed(_io_rd_big_0_T_45); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_23 = big_typ ? $signed(_io_rd_big_1_T_47) : $signed(_io_rd_big_0_T_47); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_24 = big_typ ? $signed(_io_rd_big_1_T_49) : $signed(_io_rd_big_0_T_49); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_25 = big_typ ? $signed(_io_rd_big_1_T_51) : $signed(_io_rd_big_0_T_51); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_26 = big_typ ? $signed(_io_rd_big_1_T_53) : $signed(_io_rd_big_0_T_53); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_27 = big_typ ? $signed(_io_rd_big_1_T_55) : $signed(_io_rd_big_0_T_55); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_28 = big_typ ? $signed(_io_rd_big_1_T_57) : $signed(_io_rd_big_0_T_57); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_29 = big_typ ? $signed(_io_rd_big_1_T_59) : $signed(_io_rd_big_0_T_59); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_30 = big_typ ? $signed(_io_rd_big_1_T_61) : $signed(_io_rd_big_0_T_61); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_31 = big_typ ? $signed(_io_rd_big_1_T_63) : $signed(_io_rd_big_0_T_63); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_32 = big_typ ? $signed(_io_rd_big_1_T_65) : $signed(_io_rd_big_0_T_65); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_33 = big_typ ? $signed(_io_rd_big_1_T_67) : $signed(_io_rd_big_0_T_67); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_34 = big_typ ? $signed(_io_rd_big_1_T_69) : $signed(_io_rd_big_0_T_69); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_35 = big_typ ? $signed(_io_rd_big_1_T_71) : $signed(_io_rd_big_0_T_71); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_36 = big_typ ? $signed(_io_rd_big_1_T_73) : $signed(_io_rd_big_0_T_73); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_37 = big_typ ? $signed(_io_rd_big_1_T_75) : $signed(_io_rd_big_0_T_75); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_38 = big_typ ? $signed(_io_rd_big_1_T_77) : $signed(_io_rd_big_0_T_77); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_39 = big_typ ? $signed(_io_rd_big_1_T_79) : $signed(_io_rd_big_0_T_79); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_40 = big_typ ? $signed(_io_rd_big_1_T_81) : $signed(_io_rd_big_0_T_81); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_41 = big_typ ? $signed(_io_rd_big_1_T_83) : $signed(_io_rd_big_0_T_83); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_42 = big_typ ? $signed(_io_rd_big_1_T_85) : $signed(_io_rd_big_0_T_85); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_43 = big_typ ? $signed(_io_rd_big_1_T_87) : $signed(_io_rd_big_0_T_87); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_44 = big_typ ? $signed(_io_rd_big_1_T_89) : $signed(_io_rd_big_0_T_89); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_45 = big_typ ? $signed(_io_rd_big_1_T_91) : $signed(_io_rd_big_0_T_91); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_46 = big_typ ? $signed(_io_rd_big_1_T_93) : $signed(_io_rd_big_0_T_93); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_big_1_data_47 = big_typ ? $signed(_io_rd_big_1_T_95) : $signed(_io_rd_big_0_T_95); // @[bram.scala 134:24 bram.scala 136:22 bram.scala 138:22]
  assign io_rd_small_0_0_data_0 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_10) : $signed(
    _io_rd_small_0_0_T_78_data_0); // @[Mux.scala 98:16]
  assign io_rd_small_0_0_data_1 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_12) : $signed(
    _io_rd_small_0_0_T_78_data_1); // @[Mux.scala 98:16]
  assign io_rd_small_0_0_data_2 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_14) : $signed(
    _io_rd_small_0_0_T_78_data_2); // @[Mux.scala 98:16]
  assign io_rd_small_0_0_data_3 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_16) : $signed(
    _io_rd_small_0_0_T_78_data_3); // @[Mux.scala 98:16]
  assign io_rd_small_0_0_data_4 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_18) : $signed(
    _io_rd_small_0_0_T_78_data_4); // @[Mux.scala 98:16]
  assign io_rd_small_0_0_data_5 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_20) : $signed(
    _io_rd_small_0_0_T_78_data_5); // @[Mux.scala 98:16]
  assign io_rd_small_0_0_data_6 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_22) : $signed(
    _io_rd_small_0_0_T_78_data_6); // @[Mux.scala 98:16]
  assign io_rd_small_0_0_data_7 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_24) : $signed(
    _io_rd_small_0_0_T_78_data_7); // @[Mux.scala 98:16]
  assign io_rd_small_0_1_data_0 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_27) : $signed(
    _io_rd_small_0_1_T_78_data_0); // @[Mux.scala 98:16]
  assign io_rd_small_0_1_data_1 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_29) : $signed(
    _io_rd_small_0_1_T_78_data_1); // @[Mux.scala 98:16]
  assign io_rd_small_0_1_data_2 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_31) : $signed(
    _io_rd_small_0_1_T_78_data_2); // @[Mux.scala 98:16]
  assign io_rd_small_0_1_data_3 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_33) : $signed(
    _io_rd_small_0_1_T_78_data_3); // @[Mux.scala 98:16]
  assign io_rd_small_0_1_data_4 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_35) : $signed(
    _io_rd_small_0_1_T_78_data_4); // @[Mux.scala 98:16]
  assign io_rd_small_0_1_data_5 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_37) : $signed(
    _io_rd_small_0_1_T_78_data_5); // @[Mux.scala 98:16]
  assign io_rd_small_0_1_data_6 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_39) : $signed(
    _io_rd_small_0_1_T_78_data_6); // @[Mux.scala 98:16]
  assign io_rd_small_0_1_data_7 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_41) : $signed(
    _io_rd_small_0_1_T_78_data_7); // @[Mux.scala 98:16]
  assign io_rd_small_0_2_data_0 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_44) : $signed(
    _io_rd_small_0_2_T_78_data_0); // @[Mux.scala 98:16]
  assign io_rd_small_0_2_data_1 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_46) : $signed(
    _io_rd_small_0_2_T_78_data_1); // @[Mux.scala 98:16]
  assign io_rd_small_0_2_data_2 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_48) : $signed(
    _io_rd_small_0_2_T_78_data_2); // @[Mux.scala 98:16]
  assign io_rd_small_0_2_data_3 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_50) : $signed(
    _io_rd_small_0_2_T_78_data_3); // @[Mux.scala 98:16]
  assign io_rd_small_0_2_data_4 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_52) : $signed(
    _io_rd_small_0_2_T_78_data_4); // @[Mux.scala 98:16]
  assign io_rd_small_0_2_data_5 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_54) : $signed(
    _io_rd_small_0_2_T_78_data_5); // @[Mux.scala 98:16]
  assign io_rd_small_0_2_data_6 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_56) : $signed(
    _io_rd_small_0_2_T_78_data_6); // @[Mux.scala 98:16]
  assign io_rd_small_0_2_data_7 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_58) : $signed(
    _io_rd_small_0_2_T_78_data_7); // @[Mux.scala 98:16]
  assign io_rd_small_0_3_data_0 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_61) : $signed(
    _io_rd_small_0_3_T_78_data_0); // @[Mux.scala 98:16]
  assign io_rd_small_0_3_data_1 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_63) : $signed(
    _io_rd_small_0_3_T_78_data_1); // @[Mux.scala 98:16]
  assign io_rd_small_0_3_data_2 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_65) : $signed(
    _io_rd_small_0_3_T_78_data_2); // @[Mux.scala 98:16]
  assign io_rd_small_0_3_data_3 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_67) : $signed(
    _io_rd_small_0_3_T_78_data_3); // @[Mux.scala 98:16]
  assign io_rd_small_0_3_data_4 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_69) : $signed(
    _io_rd_small_0_3_T_78_data_4); // @[Mux.scala 98:16]
  assign io_rd_small_0_3_data_5 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_71) : $signed(
    _io_rd_small_0_3_T_78_data_5); // @[Mux.scala 98:16]
  assign io_rd_small_0_3_data_6 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_73) : $signed(
    _io_rd_small_0_3_T_78_data_6); // @[Mux.scala 98:16]
  assign io_rd_small_0_3_data_7 = _io_rd_small_0_0_T_8 ? $signed(_io_rd_small_0_0_T_75) : $signed(
    _io_rd_small_0_3_T_78_data_7); // @[Mux.scala 98:16]
  assign io_rd_small_1_0_data_0 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_10) : $signed(
    _io_rd_small_1_0_T_78_data_0); // @[Mux.scala 98:16]
  assign io_rd_small_1_0_data_1 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_12) : $signed(
    _io_rd_small_1_0_T_78_data_1); // @[Mux.scala 98:16]
  assign io_rd_small_1_0_data_2 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_14) : $signed(
    _io_rd_small_1_0_T_78_data_2); // @[Mux.scala 98:16]
  assign io_rd_small_1_0_data_3 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_16) : $signed(
    _io_rd_small_1_0_T_78_data_3); // @[Mux.scala 98:16]
  assign io_rd_small_1_0_data_4 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_18) : $signed(
    _io_rd_small_1_0_T_78_data_4); // @[Mux.scala 98:16]
  assign io_rd_small_1_0_data_5 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_20) : $signed(
    _io_rd_small_1_0_T_78_data_5); // @[Mux.scala 98:16]
  assign io_rd_small_1_0_data_6 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_22) : $signed(
    _io_rd_small_1_0_T_78_data_6); // @[Mux.scala 98:16]
  assign io_rd_small_1_0_data_7 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_24) : $signed(
    _io_rd_small_1_0_T_78_data_7); // @[Mux.scala 98:16]
  assign io_rd_small_1_1_data_0 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_27) : $signed(
    _io_rd_small_1_1_T_78_data_0); // @[Mux.scala 98:16]
  assign io_rd_small_1_1_data_1 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_29) : $signed(
    _io_rd_small_1_1_T_78_data_1); // @[Mux.scala 98:16]
  assign io_rd_small_1_1_data_2 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_31) : $signed(
    _io_rd_small_1_1_T_78_data_2); // @[Mux.scala 98:16]
  assign io_rd_small_1_1_data_3 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_33) : $signed(
    _io_rd_small_1_1_T_78_data_3); // @[Mux.scala 98:16]
  assign io_rd_small_1_1_data_4 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_35) : $signed(
    _io_rd_small_1_1_T_78_data_4); // @[Mux.scala 98:16]
  assign io_rd_small_1_1_data_5 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_37) : $signed(
    _io_rd_small_1_1_T_78_data_5); // @[Mux.scala 98:16]
  assign io_rd_small_1_1_data_6 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_39) : $signed(
    _io_rd_small_1_1_T_78_data_6); // @[Mux.scala 98:16]
  assign io_rd_small_1_1_data_7 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_41) : $signed(
    _io_rd_small_1_1_T_78_data_7); // @[Mux.scala 98:16]
  assign io_rd_small_1_2_data_0 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_44) : $signed(
    _io_rd_small_1_2_T_78_data_0); // @[Mux.scala 98:16]
  assign io_rd_small_1_2_data_1 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_46) : $signed(
    _io_rd_small_1_2_T_78_data_1); // @[Mux.scala 98:16]
  assign io_rd_small_1_2_data_2 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_48) : $signed(
    _io_rd_small_1_2_T_78_data_2); // @[Mux.scala 98:16]
  assign io_rd_small_1_2_data_3 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_50) : $signed(
    _io_rd_small_1_2_T_78_data_3); // @[Mux.scala 98:16]
  assign io_rd_small_1_2_data_4 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_52) : $signed(
    _io_rd_small_1_2_T_78_data_4); // @[Mux.scala 98:16]
  assign io_rd_small_1_2_data_5 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_54) : $signed(
    _io_rd_small_1_2_T_78_data_5); // @[Mux.scala 98:16]
  assign io_rd_small_1_2_data_6 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_56) : $signed(
    _io_rd_small_1_2_T_78_data_6); // @[Mux.scala 98:16]
  assign io_rd_small_1_2_data_7 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_58) : $signed(
    _io_rd_small_1_2_T_78_data_7); // @[Mux.scala 98:16]
  assign io_rd_small_1_3_data_0 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_61) : $signed(
    _io_rd_small_1_3_T_78_data_0); // @[Mux.scala 98:16]
  assign io_rd_small_1_3_data_1 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_63) : $signed(
    _io_rd_small_1_3_T_78_data_1); // @[Mux.scala 98:16]
  assign io_rd_small_1_3_data_2 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_65) : $signed(
    _io_rd_small_1_3_T_78_data_2); // @[Mux.scala 98:16]
  assign io_rd_small_1_3_data_3 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_67) : $signed(
    _io_rd_small_1_3_T_78_data_3); // @[Mux.scala 98:16]
  assign io_rd_small_1_3_data_4 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_69) : $signed(
    _io_rd_small_1_3_T_78_data_4); // @[Mux.scala 98:16]
  assign io_rd_small_1_3_data_5 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_71) : $signed(
    _io_rd_small_1_3_T_78_data_5); // @[Mux.scala 98:16]
  assign io_rd_small_1_3_data_6 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_73) : $signed(
    _io_rd_small_1_3_T_78_data_6); // @[Mux.scala 98:16]
  assign io_rd_small_1_3_data_7 = _io_rd_small_1_0_T_8 ? $signed(_io_rd_small_1_0_T_75) : $signed(
    _io_rd_small_1_3_T_78_data_7); // @[Mux.scala 98:16]
  assign bram_big_bank0_addra = 10'h0;
  assign bram_big_bank0_clka = 1'h0;
  assign bram_big_bank0_dina = 768'h0;
  assign bram_big_bank0_wea = 1'h0;
  assign bram_big_bank0_addrb = 10'h0;
  assign bram_big_bank0_clkb = 1'h0;
  assign bram_big_bank0_dinb = 768'h0;
  assign bram_big_bank0_web = 1'h0;
  assign bram_big_bank0_1_addra = 10'h0;
  assign bram_big_bank0_1_clka = 1'h0;
  assign bram_big_bank0_1_dina = 768'h0;
  assign bram_big_bank0_1_wea = 1'h0;
  assign bram_big_bank0_1_addrb = 10'h0;
  assign bram_big_bank0_1_clkb = 1'h0;
  assign bram_big_bank0_1_dinb = 768'h0;
  assign bram_big_bank0_1_web = 1'h0;
  assign bram_small_bank0_addra = 9'h0;
  assign bram_small_bank0_clka = 1'h0;
  assign bram_small_bank0_dina = 128'h0;
  assign bram_small_bank0_wea = 1'h0;
  assign bram_small_bank0_addrb = 9'h0;
  assign bram_small_bank0_clkb = 1'h0;
  assign bram_small_bank0_dinb = 128'h0;
  assign bram_small_bank0_web = 1'h0;
  assign bram_small_bank1_addra = 9'h0;
  assign bram_small_bank1_clka = 1'h0;
  assign bram_small_bank1_dina = 128'h0;
  assign bram_small_bank1_wea = 1'h0;
  assign bram_small_bank1_addrb = 9'h0;
  assign bram_small_bank1_clkb = 1'h0;
  assign bram_small_bank1_dinb = 128'h0;
  assign bram_small_bank1_web = 1'h0;
  assign bram_small_bank2_addra = 9'h0;
  assign bram_small_bank2_clka = 1'h0;
  assign bram_small_bank2_dina = 128'h0;
  assign bram_small_bank2_wea = 1'h0;
  assign bram_small_bank2_addrb = 9'h0;
  assign bram_small_bank2_clkb = 1'h0;
  assign bram_small_bank2_dinb = 128'h0;
  assign bram_small_bank2_web = 1'h0;
  assign bram_small_bank3_addra = 9'h0;
  assign bram_small_bank3_clka = 1'h0;
  assign bram_small_bank3_dina = 128'h0;
  assign bram_small_bank3_wea = 1'h0;
  assign bram_small_bank3_addrb = 9'h0;
  assign bram_small_bank3_clkb = 1'h0;
  assign bram_small_bank3_dinb = 128'h0;
  assign bram_small_bank3_web = 1'h0;
  assign bram_small_bank4_addra = 9'h0;
  assign bram_small_bank4_clka = 1'h0;
  assign bram_small_bank4_dina = 128'h0;
  assign bram_small_bank4_wea = 1'h0;
  assign bram_small_bank4_addrb = 9'h0;
  assign bram_small_bank4_clkb = 1'h0;
  assign bram_small_bank4_dinb = 128'h0;
  assign bram_small_bank4_web = 1'h0;
  assign bram_small_bank5_addra = 9'h0;
  assign bram_small_bank5_clka = 1'h0;
  assign bram_small_bank5_dina = 128'h0;
  assign bram_small_bank5_wea = 1'h0;
  assign bram_small_bank5_addrb = 9'h0;
  assign bram_small_bank5_clkb = 1'h0;
  assign bram_small_bank5_dinb = 128'h0;
  assign bram_small_bank5_web = 1'h0;
  assign bram_small_bank6_addra = 9'h0;
  assign bram_small_bank6_clka = 1'h0;
  assign bram_small_bank6_dina = 128'h0;
  assign bram_small_bank6_wea = 1'h0;
  assign bram_small_bank6_addrb = 9'h0;
  assign bram_small_bank6_clkb = 1'h0;
  assign bram_small_bank6_dinb = 128'h0;
  assign bram_small_bank6_web = 1'h0;
  assign bram_small_bank7_addra = 9'h0;
  assign bram_small_bank7_clka = 1'h0;
  assign bram_small_bank7_dina = 128'h0;
  assign bram_small_bank7_wea = 1'h0;
  assign bram_small_bank7_addrb = 9'h0;
  assign bram_small_bank7_clkb = 1'h0;
  assign bram_small_bank7_dinb = 128'h0;
  assign bram_small_bank7_web = 1'h0;
  always @(posedge clock) begin
    if (reset) begin // @[bram.scala 87:28]
      reg_valid <= 1'h0; // @[bram.scala 87:28]
    end else begin
      reg_valid <= io_rd_valid_in; // @[bram.scala 87:28]
    end
    if (reset) begin // @[bram.scala 122:26]
      big_typ <= 1'h0; // @[bram.scala 122:26]
    end else begin
      big_typ <= _T_160;
    end
    if (reset) begin // @[bram.scala 143:22]
      typ_0 <= 2'h0; // @[bram.scala 143:22]
    end else begin
      typ_0 <= io_rd_addr1_addrs_1_addr[1:0]; // @[bram.scala 144:12]
    end
    if (reset) begin // @[bram.scala 143:22]
      typ_1 <= 2'h0; // @[bram.scala 143:22]
    end else begin
      typ_1 <= io_rd_addr2_addrs_1_addr[1:0]; // @[bram.scala 145:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  big_typ = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  typ_0 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  typ_1 = _RAND_3[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input   clock,
  input   reset,
  output  io_complete
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  GraphReader_clock; // @[top.scala 14:25]
  wire  GraphReader_reset; // @[top.scala 14:25]
  wire  GraphReader_io_valid_in; // @[top.scala 14:25]
  wire  GraphReader_io_valid_out; // @[top.scala 14:25]
  wire  GraphReader_io_flag_job; // @[top.scala 14:25]
  wire [2:0] GraphReader_io_job_big_bank_id; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_big_cnt_x_end; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_big_cnt_y_end; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_big_cnt_ic_end; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_big_cnt_loop_end; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_big_begin_loop; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_small_0_max_addr; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_small_0_cnt_y_end; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_small_0_cnt_ic_end; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_small_0_cnt_loop_end; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_small_0_begin_loop; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_job_small_0_cnt_invalid_end; // @[top.scala 14:25]
  wire [2:0] GraphReader_io_to_banks_addrs_0_bank_id; // @[top.scala 14:25]
  wire [9:0] GraphReader_io_to_banks_addrs_1_addr; // @[top.scala 14:25]
  wire  GraphReader_1_clock; // @[top.scala 15:25]
  wire  GraphReader_1_reset; // @[top.scala 15:25]
  wire  GraphReader_1_io_valid_in; // @[top.scala 15:25]
  wire  GraphReader_1_io_valid_out; // @[top.scala 15:25]
  wire  GraphReader_1_io_flag_job; // @[top.scala 15:25]
  wire [2:0] GraphReader_1_io_job_big_bank_id; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_big_cnt_x_end; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_big_cnt_y_end; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_big_cnt_ic_end; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_big_cnt_loop_end; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_big_begin_loop; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_small_0_max_addr; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_small_0_cnt_y_end; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_small_0_cnt_ic_end; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_small_0_cnt_loop_end; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_small_0_begin_loop; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_job_small_0_cnt_invalid_end; // @[top.scala 15:25]
  wire [2:0] GraphReader_1_io_to_banks_addrs_0_bank_id; // @[top.scala 15:25]
  wire [9:0] GraphReader_1_io_to_banks_addrs_1_addr; // @[top.scala 15:25]
  wire  PackReadData_clock; // @[top.scala 16:27]
  wire  PackReadData_reset; // @[top.scala 16:27]
  wire  PackReadData_io_valid_in; // @[top.scala 16:27]
  wire  PackReadData_io_valid_out; // @[top.scala 16:27]
  wire  PackReadData_io_flag_job; // @[top.scala 16:27]
  wire [9:0] PackReadData_io_job_cnt_x_end; // @[top.scala 16:27]
  wire [9:0] PackReadData_io_job_cnt_y_end; // @[top.scala 16:27]
  wire [9:0] PackReadData_io_job_in_chan; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_8; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_9; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_10; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_11; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_12; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_13; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_14; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_15; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_16; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_17; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_18; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_19; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_20; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_21; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_22; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_23; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_24; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_25; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_26; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_27; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_28; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_29; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_30; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_31; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_32; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_33; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_34; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_35; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_36; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_37; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_38; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_39; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_40; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_41; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_42; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_43; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_44; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_45; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_46; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_0_data_47; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_8; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_9; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_10; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_11; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_12; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_13; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_14; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_15; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_16; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_17; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_18; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_19; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_20; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_21; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_22; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_23; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_24; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_25; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_26; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_27; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_28; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_29; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_30; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_31; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_32; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_33; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_34; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_35; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_36; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_37; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_38; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_39; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_40; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_41; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_42; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_43; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_44; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_45; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_46; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_big_1_data_47; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_0_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_0_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_0_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_0_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_0_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_0_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_0_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_0_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_1_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_1_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_1_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_1_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_1_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_1_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_1_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_1_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_2_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_2_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_2_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_2_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_2_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_2_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_2_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_2_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_3_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_3_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_3_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_3_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_3_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_3_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_3_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_0_3_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_0_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_0_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_0_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_0_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_0_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_0_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_0_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_0_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_1_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_1_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_1_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_1_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_1_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_1_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_1_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_1_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_2_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_2_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_2_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_2_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_2_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_2_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_2_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_2_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_3_data_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_3_data_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_3_data_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_3_data_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_3_data_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_3_data_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_3_data_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_from_small_1_3_data_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_8; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_9; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_10; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_11; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_12; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_13; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_14; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_15; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_16; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_17; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_18; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_19; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_20; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_21; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_22; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_23; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_24; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_25; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_26; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_27; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_28; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_29; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_30; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_31; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_32; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_33; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_34; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_35; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_36; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_37; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_38; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_39; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_40; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_41; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_42; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_43; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_44; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_45; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_46; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_47; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_48; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_49; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_50; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_51; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_52; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_53; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_54; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_55; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_56; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_57; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_58; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_59; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_60; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_61; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_62; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_mat_63; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_8; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_up_9; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_8; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_down_9; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_left_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_left_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_left_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_left_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_left_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_left_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_left_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_left_7; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_right_0; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_right_1; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_right_2; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_right_3; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_right_4; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_right_5; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_right_6; // @[top.scala 16:27]
  wire [15:0] PackReadData_io_output_right_7; // @[top.scala 16:27]
  wire  ReadSwitch_clock; // @[top.scala 17:29]
  wire  ReadSwitch_reset; // @[top.scala 17:29]
  wire  ReadSwitch_io_flag_job; // @[top.scala 17:29]
  wire [1:0] ReadSwitch_io_job; // @[top.scala 17:29]
  wire  ReadSwitch_io_valid_in; // @[top.scala 17:29]
  wire  ReadSwitch_io_valid_out_calc8x8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_10; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_11; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_12; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_13; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_14; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_15; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_16; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_17; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_18; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_19; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_20; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_21; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_22; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_23; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_24; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_25; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_26; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_27; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_28; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_29; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_30; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_31; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_32; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_33; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_34; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_35; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_36; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_37; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_38; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_39; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_40; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_41; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_42; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_43; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_44; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_45; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_46; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_47; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_48; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_49; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_50; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_51; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_52; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_53; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_54; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_55; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_56; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_57; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_58; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_59; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_60; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_61; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_62; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_mat_63; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_up_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_down_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_left_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_left_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_left_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_left_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_left_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_left_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_left_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_left_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_right_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_right_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_right_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_right_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_right_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_right_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_right_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_right_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_from_weight_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_10; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_11; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_12; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_13; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_14; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_15; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_16; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_17; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_18; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_19; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_20; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_21; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_22; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_23; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_24; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_25; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_26; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_27; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_28; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_29; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_30; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_31; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_32; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_33; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_34; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_35; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_36; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_37; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_38; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_39; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_40; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_41; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_42; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_43; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_44; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_45; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_46; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_47; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_48; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_49; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_50; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_51; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_52; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_53; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_54; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_55; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_56; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_57; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_58; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_59; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_60; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_61; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_62; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_mat_63; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_up_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_down_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_left_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_left_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_left_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_left_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_left_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_left_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_left_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_left_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_right_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_right_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_right_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_right_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_right_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_right_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_right_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_calc8x8_right_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_10; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_11; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_12; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_13; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_14; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_0_real_15; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_10; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_11; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_12; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_13; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_14; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_1_real_15; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_10; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_11; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_12; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_13; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_14; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_2_real_15; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_0; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_1; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_2; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_3; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_4; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_5; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_6; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_7; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_8; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_9; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_10; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_11; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_12; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_13; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_14; // @[top.scala 17:29]
  wire [15:0] ReadSwitch_io_to_weight_3_real_15; // @[top.scala 17:29]
  wire  WeightReader_clock; // @[top.scala 18:29]
  wire  WeightReader_reset; // @[top.scala 18:29]
  wire  WeightReader_io_valid_in; // @[top.scala 18:29]
  wire  WeightReader_io_flag_job; // @[top.scala 18:29]
  wire [13:0] WeightReader_io_addr_end; // @[top.scala 18:29]
  wire [13:0] WeightReader_io_addr; // @[top.scala 18:29]
  wire  Calc8x8_clock; // @[top.scala 19:25]
  wire  Calc8x8_reset; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_7; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_8; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_9; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_10; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_11; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_12; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_13; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_14; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_15; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_16; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_17; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_18; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_19; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_20; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_21; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_22; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_23; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_24; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_25; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_26; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_27; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_28; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_29; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_30; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_31; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_32; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_33; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_34; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_35; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_36; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_37; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_38; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_39; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_40; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_41; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_42; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_43; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_44; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_45; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_46; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_47; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_48; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_49; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_50; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_51; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_52; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_53; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_54; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_55; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_56; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_57; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_58; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_59; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_60; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_61; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_62; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_mat_63; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_7; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_8; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_up_9; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_7; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_8; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_down_9; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_left_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_left_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_left_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_left_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_left_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_left_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_left_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_left_7; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_right_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_right_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_right_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_right_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_right_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_right_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_right_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_input_right_7; // @[top.scala 19:25]
  wire [1:0] Calc8x8_io_flag; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_7; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_8; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_9; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_10; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_11; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_12; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_13; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_14; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_0_real_15; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_7; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_8; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_9; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_10; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_11; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_12; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_13; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_14; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_1_real_15; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_7; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_8; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_9; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_10; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_11; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_12; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_13; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_14; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_2_real_15; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_0; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_1; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_2; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_3; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_4; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_5; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_6; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_7; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_8; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_9; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_10; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_11; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_12; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_13; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_14; // @[top.scala 19:25]
  wire [15:0] Calc8x8_io_weight_3_real_15; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_0; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_1; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_2; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_3; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_4; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_5; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_6; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_7; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_8; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_9; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_10; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_11; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_12; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_13; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_14; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_15; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_16; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_17; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_18; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_19; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_20; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_21; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_22; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_23; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_24; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_25; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_26; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_27; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_28; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_29; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_30; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_31; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_32; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_33; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_34; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_35; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_36; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_37; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_38; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_39; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_40; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_41; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_42; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_43; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_44; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_45; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_46; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_47; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_48; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_49; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_50; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_51; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_52; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_53; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_54; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_55; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_56; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_57; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_58; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_59; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_60; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_61; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_62; // @[top.scala 19:25]
  wire [36:0] Calc8x8_io_output_mat_63; // @[top.scala 19:25]
  wire  Calc8x8_io_valid_in; // @[top.scala 19:25]
  wire  Calc8x8_io_valid_out; // @[top.scala 19:25]
  wire  Accumu_clock; // @[top.scala 20:22]
  wire  Accumu_reset; // @[top.scala 20:22]
  wire  Accumu_io_valid_in; // @[top.scala 20:22]
  wire  Accumu_io_valid_out; // @[top.scala 20:22]
  wire  Accumu_io_flag_job; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_0; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_1; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_2; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_3; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_4; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_5; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_6; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_7; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_8; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_9; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_10; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_11; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_12; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_13; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_14; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_15; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_16; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_17; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_18; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_19; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_20; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_21; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_22; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_23; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_24; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_25; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_26; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_27; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_28; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_29; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_30; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_31; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_32; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_33; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_34; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_35; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_36; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_37; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_38; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_39; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_40; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_41; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_42; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_43; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_44; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_45; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_46; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_47; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_48; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_49; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_50; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_51; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_52; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_53; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_54; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_55; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_56; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_57; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_58; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_59; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_60; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_61; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_62; // @[top.scala 20:22]
  wire [36:0] Accumu_io_in_from_calc8x8_mat_63; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_0; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_1; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_2; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_3; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_4; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_5; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_6; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_7; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_8; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_9; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_10; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_11; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_12; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_13; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_14; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_15; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_16; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_17; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_18; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_19; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_20; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_21; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_22; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_23; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_24; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_25; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_26; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_27; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_28; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_29; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_30; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_31; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_32; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_33; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_34; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_35; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_36; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_37; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_38; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_39; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_40; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_41; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_42; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_43; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_44; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_45; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_46; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_47; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_48; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_49; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_50; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_51; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_52; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_53; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_54; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_55; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_56; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_57; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_58; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_59; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_60; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_61; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_62; // @[top.scala 20:22]
  wire [43:0] Accumu_io_result_mat_63; // @[top.scala 20:22]
  wire [9:0] Accumu_io_csum; // @[top.scala 20:22]
  wire [9:0] Accumu_io_bias_end_addr; // @[top.scala 20:22]
  wire [9:0] Accumu_io_bias_addr; // @[top.scala 20:22]
  wire [35:0] Accumu_io_bias_in; // @[top.scala 20:22]
  wire  Accumu_io_is_in_use; // @[top.scala 20:22]
  wire  Quant_clock; // @[top.scala 21:23]
  wire  Quant_reset; // @[top.scala 21:23]
  wire  Quant_io_valid_in; // @[top.scala 21:23]
  wire  Quant_io_valid_out; // @[top.scala 21:23]
  wire  Quant_io_flag_job; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_0; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_1; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_2; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_3; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_4; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_5; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_6; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_7; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_8; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_9; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_10; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_11; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_12; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_13; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_14; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_15; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_16; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_17; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_18; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_19; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_20; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_21; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_22; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_23; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_24; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_25; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_26; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_27; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_28; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_29; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_30; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_31; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_32; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_33; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_34; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_35; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_36; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_37; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_38; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_39; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_40; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_41; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_42; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_43; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_44; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_45; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_46; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_47; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_48; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_49; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_50; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_51; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_52; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_53; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_54; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_55; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_56; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_57; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_58; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_59; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_60; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_61; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_62; // @[top.scala 21:23]
  wire [43:0] Quant_io_in_from_accumu_mat_63; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_0; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_1; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_2; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_3; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_4; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_5; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_6; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_7; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_8; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_9; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_10; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_11; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_12; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_13; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_14; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_15; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_16; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_17; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_18; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_19; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_20; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_21; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_22; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_23; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_24; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_25; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_26; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_27; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_28; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_29; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_30; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_31; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_32; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_33; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_34; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_35; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_36; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_37; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_38; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_39; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_40; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_41; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_42; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_43; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_44; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_45; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_46; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_47; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_48; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_49; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_50; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_51; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_52; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_53; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_54; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_55; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_56; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_57; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_58; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_59; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_60; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_61; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_62; // @[top.scala 21:23]
  wire [15:0] Quant_io_result_mat_63; // @[top.scala 21:23]
  wire [5:0] Quant_io_quant_in_in_q; // @[top.scala 21:23]
  wire [5:0] Quant_io_quant_in_out_q; // @[top.scala 21:23]
  wire  WriteSwitch_io_valid_in_0; // @[top.scala 22:30]
  wire  WriteSwitch_io_valid_out; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_0; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_1; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_2; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_3; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_4; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_5; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_6; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_7; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_8; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_9; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_10; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_11; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_12; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_13; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_14; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_15; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_16; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_17; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_18; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_19; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_20; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_21; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_22; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_23; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_24; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_25; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_26; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_27; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_28; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_29; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_30; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_31; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_32; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_33; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_34; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_35; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_36; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_37; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_38; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_39; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_40; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_41; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_42; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_43; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_44; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_45; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_46; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_47; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_48; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_49; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_50; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_51; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_52; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_53; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_54; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_55; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_56; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_57; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_58; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_59; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_60; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_61; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_62; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_input_0_mat_63; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_0; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_1; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_2; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_3; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_4; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_5; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_6; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_7; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_8; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_9; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_10; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_11; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_12; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_13; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_14; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_15; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_16; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_17; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_18; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_19; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_20; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_21; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_22; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_23; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_24; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_25; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_26; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_27; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_28; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_29; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_30; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_31; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_32; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_33; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_34; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_35; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_36; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_37; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_38; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_39; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_40; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_41; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_42; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_43; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_44; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_45; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_46; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_47; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_48; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_49; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_50; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_51; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_52; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_53; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_54; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_55; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_56; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_57; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_58; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_59; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_60; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_61; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_62; // @[top.scala 22:30]
  wire [15:0] WriteSwitch_io_output_mat_63; // @[top.scala 22:30]
  wire  RealWriter_clock; // @[top.scala 23:24]
  wire  RealWriter_reset; // @[top.scala 23:24]
  wire  RealWriter_io_valid_in; // @[top.scala 23:24]
  wire  RealWriter_io_valid_out; // @[top.scala 23:24]
  wire  RealWriter_io_flag_job; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_0; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_1; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_2; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_3; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_4; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_5; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_6; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_7; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_8; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_9; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_10; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_11; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_12; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_13; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_14; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_15; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_16; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_17; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_18; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_19; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_20; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_21; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_22; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_23; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_24; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_25; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_26; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_27; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_28; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_29; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_30; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_31; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_32; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_33; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_34; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_35; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_36; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_37; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_38; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_39; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_40; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_41; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_42; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_43; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_44; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_45; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_46; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_47; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_48; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_49; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_50; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_51; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_52; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_53; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_54; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_55; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_56; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_57; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_58; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_59; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_60; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_61; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_62; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_in_from_quant_mat_63; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_big_begin_addr; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_big_max_addr; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_big_cnt_ic_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_big_a; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_0_begin_addr; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_0_max_addr; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_0_cnt_y_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_0_cnt_ic_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_0_a; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_job_job_0_small_0_ano_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_1_begin_addr; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_1_max_addr; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_job_job_0_small_1_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_1_cnt_y_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_1_cnt_ic_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_0_small_1_a; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_job_job_0_small_1_ano_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_big_begin_addr; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_big_max_addr; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_job_job_1_big_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_big_cnt_ic_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_big_a; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_0_begin_addr; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_0_max_addr; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_job_job_1_small_0_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_0_cnt_y_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_0_cnt_ic_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_0_a; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_job_job_1_small_0_ano_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_1_begin_addr; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_1_max_addr; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_job_job_1_small_1_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_1_cnt_y_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_1_cnt_ic_end; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_job_1_small_1_a; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_job_job_1_small_1_ano_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_job_out_chan; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_0; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_1; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_2; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_3; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_4; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_5; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_6; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_7; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_8; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_9; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_10; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_11; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_12; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_13; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_14; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_15; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_16; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_17; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_18; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_19; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_20; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_21; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_22; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_23; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_24; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_25; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_26; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_27; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_28; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_29; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_30; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_31; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_32; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_33; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_34; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_35; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_36; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_37; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_38; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_39; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_40; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_41; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_42; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_43; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_44; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_45; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_46; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_bigbank_data_47; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_0_data_0; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_0_data_1; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_0_data_2; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_0_data_3; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_0_data_4; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_0_data_5; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_0_data_6; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_0_data_7; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_1_data_0; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_1_data_1; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_1_data_2; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_1_data_3; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_1_data_4; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_1_data_5; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_1_data_6; // @[top.scala 23:24]
  wire [15:0] RealWriter_io_to_smallbank_1_data_7; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_to_banks_addrs_0_addr; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_to_banks_addrs_0_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_to_banks_addrs_1_addr; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_to_banks_addrs_1_bank_id; // @[top.scala 23:24]
  wire [9:0] RealWriter_io_to_banks_addrs_2_addr; // @[top.scala 23:24]
  wire [2:0] RealWriter_io_to_banks_addrs_2_bank_id; // @[top.scala 23:24]
  wire  ROMWeight_clock; // @[top.scala 26:28]
  wire [13:0] ROMWeight_io_addr; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_0; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_1; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_2; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_3; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_4; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_5; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_6; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_7; // @[top.scala 26:28]
  wire [15:0] ROMWeight_io_out_8; // @[top.scala 26:28]
  wire  ROMBias_clock; // @[top.scala 27:26]
  wire [7:0] ROMBias_io_addr; // @[top.scala 27:26]
  wire [35:0] ROMBias_io_out; // @[top.scala 27:26]
  wire  RAMGroup_clock; // @[top.scala 28:22]
  wire  RAMGroup_reset; // @[top.scala 28:22]
  wire  RAMGroup_io_rd_valid_in; // @[top.scala 28:22]
  wire  RAMGroup_io_rd_valid_out; // @[top.scala 28:22]
  wire [2:0] RAMGroup_io_rd_addr1_addrs_0_bank_id; // @[top.scala 28:22]
  wire [9:0] RAMGroup_io_rd_addr1_addrs_1_addr; // @[top.scala 28:22]
  wire [9:0] RAMGroup_io_rd_addr2_addrs_1_addr; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_8; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_9; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_10; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_11; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_12; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_13; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_14; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_15; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_16; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_17; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_18; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_19; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_20; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_21; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_22; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_23; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_24; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_25; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_26; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_27; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_28; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_29; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_30; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_31; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_32; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_33; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_34; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_35; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_36; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_37; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_38; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_39; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_40; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_41; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_42; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_43; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_44; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_45; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_46; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_0_data_47; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_8; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_9; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_10; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_11; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_12; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_13; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_14; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_15; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_16; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_17; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_18; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_19; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_20; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_21; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_22; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_23; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_24; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_25; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_26; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_27; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_28; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_29; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_30; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_31; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_32; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_33; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_34; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_35; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_36; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_37; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_38; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_39; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_40; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_41; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_42; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_43; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_44; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_45; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_46; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_big_1_data_47; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_0_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_0_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_0_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_0_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_0_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_0_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_0_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_0_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_1_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_1_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_1_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_1_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_1_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_1_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_1_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_1_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_2_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_2_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_2_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_2_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_2_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_2_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_2_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_2_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_3_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_3_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_3_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_3_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_3_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_3_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_3_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_0_3_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_0_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_0_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_0_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_0_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_0_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_0_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_0_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_0_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_1_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_1_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_1_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_1_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_1_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_1_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_1_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_1_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_2_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_2_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_2_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_2_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_2_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_2_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_2_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_2_data_7; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_3_data_0; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_3_data_1; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_3_data_2; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_3_data_3; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_3_data_4; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_3_data_5; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_3_data_6; // @[top.scala 28:22]
  wire [15:0] RAMGroup_io_rd_small_1_3_data_7; // @[top.scala 28:22]
  reg [9:0] counter_ccnt; // @[top.scala 134:26]
  reg [9:0] counter_cend; // @[top.scala 134:26]
  reg [2:0] state; // @[top.scala 135:24]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  nxt = counter_ccnt == counter_cend; // @[utils.scala 17:20]
  wire [9:0] _counter_ccnt_T_1 = counter_ccnt + 10'h1; // @[utils.scala 18:35]
  wire [9:0] _counter_ccnt_T_2 = nxt ? 10'h0 : _counter_ccnt_T_1; // @[utils.scala 18:20]
  wire [2:0] _GEN_0 = nxt ? 3'h2 : state; // @[top.scala 153:36 top.scala 155:27 top.scala 135:24]
  wire  _T_2 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_7 = _T_1 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 top.scala 161:26 top.scala 64:18]
  wire [5:0] _GEN_148 = _T ? 6'h3f : 6'h0; // @[Conditional.scala 40:58 para.scala 74:21 top.scala 45:26]
  wire [3:0] _GEN_152 = _T ? 4'hf : 4'h0; // @[Conditional.scala 40:58 para.scala 92:17 top.scala 72:15]
  GraphReader GraphReader ( // @[top.scala 14:25]
    .clock(GraphReader_clock),
    .reset(GraphReader_reset),
    .io_valid_in(GraphReader_io_valid_in),
    .io_valid_out(GraphReader_io_valid_out),
    .io_flag_job(GraphReader_io_flag_job),
    .io_job_big_bank_id(GraphReader_io_job_big_bank_id),
    .io_job_big_cnt_x_end(GraphReader_io_job_big_cnt_x_end),
    .io_job_big_cnt_y_end(GraphReader_io_job_big_cnt_y_end),
    .io_job_big_cnt_ic_end(GraphReader_io_job_big_cnt_ic_end),
    .io_job_big_cnt_loop_end(GraphReader_io_job_big_cnt_loop_end),
    .io_job_big_begin_loop(GraphReader_io_job_big_begin_loop),
    .io_job_small_0_max_addr(GraphReader_io_job_small_0_max_addr),
    .io_job_small_0_cnt_y_end(GraphReader_io_job_small_0_cnt_y_end),
    .io_job_small_0_cnt_ic_end(GraphReader_io_job_small_0_cnt_ic_end),
    .io_job_small_0_cnt_loop_end(GraphReader_io_job_small_0_cnt_loop_end),
    .io_job_small_0_begin_loop(GraphReader_io_job_small_0_begin_loop),
    .io_job_small_0_cnt_invalid_end(GraphReader_io_job_small_0_cnt_invalid_end),
    .io_to_banks_addrs_0_bank_id(GraphReader_io_to_banks_addrs_0_bank_id),
    .io_to_banks_addrs_1_addr(GraphReader_io_to_banks_addrs_1_addr)
  );
  GraphReader GraphReader_1 ( // @[top.scala 15:25]
    .clock(GraphReader_1_clock),
    .reset(GraphReader_1_reset),
    .io_valid_in(GraphReader_1_io_valid_in),
    .io_valid_out(GraphReader_1_io_valid_out),
    .io_flag_job(GraphReader_1_io_flag_job),
    .io_job_big_bank_id(GraphReader_1_io_job_big_bank_id),
    .io_job_big_cnt_x_end(GraphReader_1_io_job_big_cnt_x_end),
    .io_job_big_cnt_y_end(GraphReader_1_io_job_big_cnt_y_end),
    .io_job_big_cnt_ic_end(GraphReader_1_io_job_big_cnt_ic_end),
    .io_job_big_cnt_loop_end(GraphReader_1_io_job_big_cnt_loop_end),
    .io_job_big_begin_loop(GraphReader_1_io_job_big_begin_loop),
    .io_job_small_0_max_addr(GraphReader_1_io_job_small_0_max_addr),
    .io_job_small_0_cnt_y_end(GraphReader_1_io_job_small_0_cnt_y_end),
    .io_job_small_0_cnt_ic_end(GraphReader_1_io_job_small_0_cnt_ic_end),
    .io_job_small_0_cnt_loop_end(GraphReader_1_io_job_small_0_cnt_loop_end),
    .io_job_small_0_begin_loop(GraphReader_1_io_job_small_0_begin_loop),
    .io_job_small_0_cnt_invalid_end(GraphReader_1_io_job_small_0_cnt_invalid_end),
    .io_to_banks_addrs_0_bank_id(GraphReader_1_io_to_banks_addrs_0_bank_id),
    .io_to_banks_addrs_1_addr(GraphReader_1_io_to_banks_addrs_1_addr)
  );
  PackReadData PackReadData ( // @[top.scala 16:27]
    .clock(PackReadData_clock),
    .reset(PackReadData_reset),
    .io_valid_in(PackReadData_io_valid_in),
    .io_valid_out(PackReadData_io_valid_out),
    .io_flag_job(PackReadData_io_flag_job),
    .io_job_cnt_x_end(PackReadData_io_job_cnt_x_end),
    .io_job_cnt_y_end(PackReadData_io_job_cnt_y_end),
    .io_job_in_chan(PackReadData_io_job_in_chan),
    .io_from_big_0_data_0(PackReadData_io_from_big_0_data_0),
    .io_from_big_0_data_1(PackReadData_io_from_big_0_data_1),
    .io_from_big_0_data_2(PackReadData_io_from_big_0_data_2),
    .io_from_big_0_data_3(PackReadData_io_from_big_0_data_3),
    .io_from_big_0_data_4(PackReadData_io_from_big_0_data_4),
    .io_from_big_0_data_5(PackReadData_io_from_big_0_data_5),
    .io_from_big_0_data_6(PackReadData_io_from_big_0_data_6),
    .io_from_big_0_data_7(PackReadData_io_from_big_0_data_7),
    .io_from_big_0_data_8(PackReadData_io_from_big_0_data_8),
    .io_from_big_0_data_9(PackReadData_io_from_big_0_data_9),
    .io_from_big_0_data_10(PackReadData_io_from_big_0_data_10),
    .io_from_big_0_data_11(PackReadData_io_from_big_0_data_11),
    .io_from_big_0_data_12(PackReadData_io_from_big_0_data_12),
    .io_from_big_0_data_13(PackReadData_io_from_big_0_data_13),
    .io_from_big_0_data_14(PackReadData_io_from_big_0_data_14),
    .io_from_big_0_data_15(PackReadData_io_from_big_0_data_15),
    .io_from_big_0_data_16(PackReadData_io_from_big_0_data_16),
    .io_from_big_0_data_17(PackReadData_io_from_big_0_data_17),
    .io_from_big_0_data_18(PackReadData_io_from_big_0_data_18),
    .io_from_big_0_data_19(PackReadData_io_from_big_0_data_19),
    .io_from_big_0_data_20(PackReadData_io_from_big_0_data_20),
    .io_from_big_0_data_21(PackReadData_io_from_big_0_data_21),
    .io_from_big_0_data_22(PackReadData_io_from_big_0_data_22),
    .io_from_big_0_data_23(PackReadData_io_from_big_0_data_23),
    .io_from_big_0_data_24(PackReadData_io_from_big_0_data_24),
    .io_from_big_0_data_25(PackReadData_io_from_big_0_data_25),
    .io_from_big_0_data_26(PackReadData_io_from_big_0_data_26),
    .io_from_big_0_data_27(PackReadData_io_from_big_0_data_27),
    .io_from_big_0_data_28(PackReadData_io_from_big_0_data_28),
    .io_from_big_0_data_29(PackReadData_io_from_big_0_data_29),
    .io_from_big_0_data_30(PackReadData_io_from_big_0_data_30),
    .io_from_big_0_data_31(PackReadData_io_from_big_0_data_31),
    .io_from_big_0_data_32(PackReadData_io_from_big_0_data_32),
    .io_from_big_0_data_33(PackReadData_io_from_big_0_data_33),
    .io_from_big_0_data_34(PackReadData_io_from_big_0_data_34),
    .io_from_big_0_data_35(PackReadData_io_from_big_0_data_35),
    .io_from_big_0_data_36(PackReadData_io_from_big_0_data_36),
    .io_from_big_0_data_37(PackReadData_io_from_big_0_data_37),
    .io_from_big_0_data_38(PackReadData_io_from_big_0_data_38),
    .io_from_big_0_data_39(PackReadData_io_from_big_0_data_39),
    .io_from_big_0_data_40(PackReadData_io_from_big_0_data_40),
    .io_from_big_0_data_41(PackReadData_io_from_big_0_data_41),
    .io_from_big_0_data_42(PackReadData_io_from_big_0_data_42),
    .io_from_big_0_data_43(PackReadData_io_from_big_0_data_43),
    .io_from_big_0_data_44(PackReadData_io_from_big_0_data_44),
    .io_from_big_0_data_45(PackReadData_io_from_big_0_data_45),
    .io_from_big_0_data_46(PackReadData_io_from_big_0_data_46),
    .io_from_big_0_data_47(PackReadData_io_from_big_0_data_47),
    .io_from_big_1_data_0(PackReadData_io_from_big_1_data_0),
    .io_from_big_1_data_1(PackReadData_io_from_big_1_data_1),
    .io_from_big_1_data_2(PackReadData_io_from_big_1_data_2),
    .io_from_big_1_data_3(PackReadData_io_from_big_1_data_3),
    .io_from_big_1_data_4(PackReadData_io_from_big_1_data_4),
    .io_from_big_1_data_5(PackReadData_io_from_big_1_data_5),
    .io_from_big_1_data_6(PackReadData_io_from_big_1_data_6),
    .io_from_big_1_data_7(PackReadData_io_from_big_1_data_7),
    .io_from_big_1_data_8(PackReadData_io_from_big_1_data_8),
    .io_from_big_1_data_9(PackReadData_io_from_big_1_data_9),
    .io_from_big_1_data_10(PackReadData_io_from_big_1_data_10),
    .io_from_big_1_data_11(PackReadData_io_from_big_1_data_11),
    .io_from_big_1_data_12(PackReadData_io_from_big_1_data_12),
    .io_from_big_1_data_13(PackReadData_io_from_big_1_data_13),
    .io_from_big_1_data_14(PackReadData_io_from_big_1_data_14),
    .io_from_big_1_data_15(PackReadData_io_from_big_1_data_15),
    .io_from_big_1_data_16(PackReadData_io_from_big_1_data_16),
    .io_from_big_1_data_17(PackReadData_io_from_big_1_data_17),
    .io_from_big_1_data_18(PackReadData_io_from_big_1_data_18),
    .io_from_big_1_data_19(PackReadData_io_from_big_1_data_19),
    .io_from_big_1_data_20(PackReadData_io_from_big_1_data_20),
    .io_from_big_1_data_21(PackReadData_io_from_big_1_data_21),
    .io_from_big_1_data_22(PackReadData_io_from_big_1_data_22),
    .io_from_big_1_data_23(PackReadData_io_from_big_1_data_23),
    .io_from_big_1_data_24(PackReadData_io_from_big_1_data_24),
    .io_from_big_1_data_25(PackReadData_io_from_big_1_data_25),
    .io_from_big_1_data_26(PackReadData_io_from_big_1_data_26),
    .io_from_big_1_data_27(PackReadData_io_from_big_1_data_27),
    .io_from_big_1_data_28(PackReadData_io_from_big_1_data_28),
    .io_from_big_1_data_29(PackReadData_io_from_big_1_data_29),
    .io_from_big_1_data_30(PackReadData_io_from_big_1_data_30),
    .io_from_big_1_data_31(PackReadData_io_from_big_1_data_31),
    .io_from_big_1_data_32(PackReadData_io_from_big_1_data_32),
    .io_from_big_1_data_33(PackReadData_io_from_big_1_data_33),
    .io_from_big_1_data_34(PackReadData_io_from_big_1_data_34),
    .io_from_big_1_data_35(PackReadData_io_from_big_1_data_35),
    .io_from_big_1_data_36(PackReadData_io_from_big_1_data_36),
    .io_from_big_1_data_37(PackReadData_io_from_big_1_data_37),
    .io_from_big_1_data_38(PackReadData_io_from_big_1_data_38),
    .io_from_big_1_data_39(PackReadData_io_from_big_1_data_39),
    .io_from_big_1_data_40(PackReadData_io_from_big_1_data_40),
    .io_from_big_1_data_41(PackReadData_io_from_big_1_data_41),
    .io_from_big_1_data_42(PackReadData_io_from_big_1_data_42),
    .io_from_big_1_data_43(PackReadData_io_from_big_1_data_43),
    .io_from_big_1_data_44(PackReadData_io_from_big_1_data_44),
    .io_from_big_1_data_45(PackReadData_io_from_big_1_data_45),
    .io_from_big_1_data_46(PackReadData_io_from_big_1_data_46),
    .io_from_big_1_data_47(PackReadData_io_from_big_1_data_47),
    .io_from_small_0_0_data_0(PackReadData_io_from_small_0_0_data_0),
    .io_from_small_0_0_data_1(PackReadData_io_from_small_0_0_data_1),
    .io_from_small_0_0_data_2(PackReadData_io_from_small_0_0_data_2),
    .io_from_small_0_0_data_3(PackReadData_io_from_small_0_0_data_3),
    .io_from_small_0_0_data_4(PackReadData_io_from_small_0_0_data_4),
    .io_from_small_0_0_data_5(PackReadData_io_from_small_0_0_data_5),
    .io_from_small_0_0_data_6(PackReadData_io_from_small_0_0_data_6),
    .io_from_small_0_0_data_7(PackReadData_io_from_small_0_0_data_7),
    .io_from_small_0_1_data_0(PackReadData_io_from_small_0_1_data_0),
    .io_from_small_0_1_data_1(PackReadData_io_from_small_0_1_data_1),
    .io_from_small_0_1_data_2(PackReadData_io_from_small_0_1_data_2),
    .io_from_small_0_1_data_3(PackReadData_io_from_small_0_1_data_3),
    .io_from_small_0_1_data_4(PackReadData_io_from_small_0_1_data_4),
    .io_from_small_0_1_data_5(PackReadData_io_from_small_0_1_data_5),
    .io_from_small_0_1_data_6(PackReadData_io_from_small_0_1_data_6),
    .io_from_small_0_1_data_7(PackReadData_io_from_small_0_1_data_7),
    .io_from_small_0_2_data_0(PackReadData_io_from_small_0_2_data_0),
    .io_from_small_0_2_data_1(PackReadData_io_from_small_0_2_data_1),
    .io_from_small_0_2_data_2(PackReadData_io_from_small_0_2_data_2),
    .io_from_small_0_2_data_3(PackReadData_io_from_small_0_2_data_3),
    .io_from_small_0_2_data_4(PackReadData_io_from_small_0_2_data_4),
    .io_from_small_0_2_data_5(PackReadData_io_from_small_0_2_data_5),
    .io_from_small_0_2_data_6(PackReadData_io_from_small_0_2_data_6),
    .io_from_small_0_2_data_7(PackReadData_io_from_small_0_2_data_7),
    .io_from_small_0_3_data_0(PackReadData_io_from_small_0_3_data_0),
    .io_from_small_0_3_data_1(PackReadData_io_from_small_0_3_data_1),
    .io_from_small_0_3_data_2(PackReadData_io_from_small_0_3_data_2),
    .io_from_small_0_3_data_3(PackReadData_io_from_small_0_3_data_3),
    .io_from_small_0_3_data_4(PackReadData_io_from_small_0_3_data_4),
    .io_from_small_0_3_data_5(PackReadData_io_from_small_0_3_data_5),
    .io_from_small_0_3_data_6(PackReadData_io_from_small_0_3_data_6),
    .io_from_small_0_3_data_7(PackReadData_io_from_small_0_3_data_7),
    .io_from_small_1_0_data_0(PackReadData_io_from_small_1_0_data_0),
    .io_from_small_1_0_data_1(PackReadData_io_from_small_1_0_data_1),
    .io_from_small_1_0_data_2(PackReadData_io_from_small_1_0_data_2),
    .io_from_small_1_0_data_3(PackReadData_io_from_small_1_0_data_3),
    .io_from_small_1_0_data_4(PackReadData_io_from_small_1_0_data_4),
    .io_from_small_1_0_data_5(PackReadData_io_from_small_1_0_data_5),
    .io_from_small_1_0_data_6(PackReadData_io_from_small_1_0_data_6),
    .io_from_small_1_0_data_7(PackReadData_io_from_small_1_0_data_7),
    .io_from_small_1_1_data_0(PackReadData_io_from_small_1_1_data_0),
    .io_from_small_1_1_data_1(PackReadData_io_from_small_1_1_data_1),
    .io_from_small_1_1_data_2(PackReadData_io_from_small_1_1_data_2),
    .io_from_small_1_1_data_3(PackReadData_io_from_small_1_1_data_3),
    .io_from_small_1_1_data_4(PackReadData_io_from_small_1_1_data_4),
    .io_from_small_1_1_data_5(PackReadData_io_from_small_1_1_data_5),
    .io_from_small_1_1_data_6(PackReadData_io_from_small_1_1_data_6),
    .io_from_small_1_1_data_7(PackReadData_io_from_small_1_1_data_7),
    .io_from_small_1_2_data_0(PackReadData_io_from_small_1_2_data_0),
    .io_from_small_1_2_data_1(PackReadData_io_from_small_1_2_data_1),
    .io_from_small_1_2_data_2(PackReadData_io_from_small_1_2_data_2),
    .io_from_small_1_2_data_3(PackReadData_io_from_small_1_2_data_3),
    .io_from_small_1_2_data_4(PackReadData_io_from_small_1_2_data_4),
    .io_from_small_1_2_data_5(PackReadData_io_from_small_1_2_data_5),
    .io_from_small_1_2_data_6(PackReadData_io_from_small_1_2_data_6),
    .io_from_small_1_2_data_7(PackReadData_io_from_small_1_2_data_7),
    .io_from_small_1_3_data_0(PackReadData_io_from_small_1_3_data_0),
    .io_from_small_1_3_data_1(PackReadData_io_from_small_1_3_data_1),
    .io_from_small_1_3_data_2(PackReadData_io_from_small_1_3_data_2),
    .io_from_small_1_3_data_3(PackReadData_io_from_small_1_3_data_3),
    .io_from_small_1_3_data_4(PackReadData_io_from_small_1_3_data_4),
    .io_from_small_1_3_data_5(PackReadData_io_from_small_1_3_data_5),
    .io_from_small_1_3_data_6(PackReadData_io_from_small_1_3_data_6),
    .io_from_small_1_3_data_7(PackReadData_io_from_small_1_3_data_7),
    .io_output_mat_0(PackReadData_io_output_mat_0),
    .io_output_mat_1(PackReadData_io_output_mat_1),
    .io_output_mat_2(PackReadData_io_output_mat_2),
    .io_output_mat_3(PackReadData_io_output_mat_3),
    .io_output_mat_4(PackReadData_io_output_mat_4),
    .io_output_mat_5(PackReadData_io_output_mat_5),
    .io_output_mat_6(PackReadData_io_output_mat_6),
    .io_output_mat_7(PackReadData_io_output_mat_7),
    .io_output_mat_8(PackReadData_io_output_mat_8),
    .io_output_mat_9(PackReadData_io_output_mat_9),
    .io_output_mat_10(PackReadData_io_output_mat_10),
    .io_output_mat_11(PackReadData_io_output_mat_11),
    .io_output_mat_12(PackReadData_io_output_mat_12),
    .io_output_mat_13(PackReadData_io_output_mat_13),
    .io_output_mat_14(PackReadData_io_output_mat_14),
    .io_output_mat_15(PackReadData_io_output_mat_15),
    .io_output_mat_16(PackReadData_io_output_mat_16),
    .io_output_mat_17(PackReadData_io_output_mat_17),
    .io_output_mat_18(PackReadData_io_output_mat_18),
    .io_output_mat_19(PackReadData_io_output_mat_19),
    .io_output_mat_20(PackReadData_io_output_mat_20),
    .io_output_mat_21(PackReadData_io_output_mat_21),
    .io_output_mat_22(PackReadData_io_output_mat_22),
    .io_output_mat_23(PackReadData_io_output_mat_23),
    .io_output_mat_24(PackReadData_io_output_mat_24),
    .io_output_mat_25(PackReadData_io_output_mat_25),
    .io_output_mat_26(PackReadData_io_output_mat_26),
    .io_output_mat_27(PackReadData_io_output_mat_27),
    .io_output_mat_28(PackReadData_io_output_mat_28),
    .io_output_mat_29(PackReadData_io_output_mat_29),
    .io_output_mat_30(PackReadData_io_output_mat_30),
    .io_output_mat_31(PackReadData_io_output_mat_31),
    .io_output_mat_32(PackReadData_io_output_mat_32),
    .io_output_mat_33(PackReadData_io_output_mat_33),
    .io_output_mat_34(PackReadData_io_output_mat_34),
    .io_output_mat_35(PackReadData_io_output_mat_35),
    .io_output_mat_36(PackReadData_io_output_mat_36),
    .io_output_mat_37(PackReadData_io_output_mat_37),
    .io_output_mat_38(PackReadData_io_output_mat_38),
    .io_output_mat_39(PackReadData_io_output_mat_39),
    .io_output_mat_40(PackReadData_io_output_mat_40),
    .io_output_mat_41(PackReadData_io_output_mat_41),
    .io_output_mat_42(PackReadData_io_output_mat_42),
    .io_output_mat_43(PackReadData_io_output_mat_43),
    .io_output_mat_44(PackReadData_io_output_mat_44),
    .io_output_mat_45(PackReadData_io_output_mat_45),
    .io_output_mat_46(PackReadData_io_output_mat_46),
    .io_output_mat_47(PackReadData_io_output_mat_47),
    .io_output_mat_48(PackReadData_io_output_mat_48),
    .io_output_mat_49(PackReadData_io_output_mat_49),
    .io_output_mat_50(PackReadData_io_output_mat_50),
    .io_output_mat_51(PackReadData_io_output_mat_51),
    .io_output_mat_52(PackReadData_io_output_mat_52),
    .io_output_mat_53(PackReadData_io_output_mat_53),
    .io_output_mat_54(PackReadData_io_output_mat_54),
    .io_output_mat_55(PackReadData_io_output_mat_55),
    .io_output_mat_56(PackReadData_io_output_mat_56),
    .io_output_mat_57(PackReadData_io_output_mat_57),
    .io_output_mat_58(PackReadData_io_output_mat_58),
    .io_output_mat_59(PackReadData_io_output_mat_59),
    .io_output_mat_60(PackReadData_io_output_mat_60),
    .io_output_mat_61(PackReadData_io_output_mat_61),
    .io_output_mat_62(PackReadData_io_output_mat_62),
    .io_output_mat_63(PackReadData_io_output_mat_63),
    .io_output_up_0(PackReadData_io_output_up_0),
    .io_output_up_1(PackReadData_io_output_up_1),
    .io_output_up_2(PackReadData_io_output_up_2),
    .io_output_up_3(PackReadData_io_output_up_3),
    .io_output_up_4(PackReadData_io_output_up_4),
    .io_output_up_5(PackReadData_io_output_up_5),
    .io_output_up_6(PackReadData_io_output_up_6),
    .io_output_up_7(PackReadData_io_output_up_7),
    .io_output_up_8(PackReadData_io_output_up_8),
    .io_output_up_9(PackReadData_io_output_up_9),
    .io_output_down_0(PackReadData_io_output_down_0),
    .io_output_down_1(PackReadData_io_output_down_1),
    .io_output_down_2(PackReadData_io_output_down_2),
    .io_output_down_3(PackReadData_io_output_down_3),
    .io_output_down_4(PackReadData_io_output_down_4),
    .io_output_down_5(PackReadData_io_output_down_5),
    .io_output_down_6(PackReadData_io_output_down_6),
    .io_output_down_7(PackReadData_io_output_down_7),
    .io_output_down_8(PackReadData_io_output_down_8),
    .io_output_down_9(PackReadData_io_output_down_9),
    .io_output_left_0(PackReadData_io_output_left_0),
    .io_output_left_1(PackReadData_io_output_left_1),
    .io_output_left_2(PackReadData_io_output_left_2),
    .io_output_left_3(PackReadData_io_output_left_3),
    .io_output_left_4(PackReadData_io_output_left_4),
    .io_output_left_5(PackReadData_io_output_left_5),
    .io_output_left_6(PackReadData_io_output_left_6),
    .io_output_left_7(PackReadData_io_output_left_7),
    .io_output_right_0(PackReadData_io_output_right_0),
    .io_output_right_1(PackReadData_io_output_right_1),
    .io_output_right_2(PackReadData_io_output_right_2),
    .io_output_right_3(PackReadData_io_output_right_3),
    .io_output_right_4(PackReadData_io_output_right_4),
    .io_output_right_5(PackReadData_io_output_right_5),
    .io_output_right_6(PackReadData_io_output_right_6),
    .io_output_right_7(PackReadData_io_output_right_7)
  );
  ReadSwitch ReadSwitch ( // @[top.scala 17:29]
    .clock(ReadSwitch_clock),
    .reset(ReadSwitch_reset),
    .io_flag_job(ReadSwitch_io_flag_job),
    .io_job(ReadSwitch_io_job),
    .io_valid_in(ReadSwitch_io_valid_in),
    .io_valid_out_calc8x8(ReadSwitch_io_valid_out_calc8x8),
    .io_from_mat_0(ReadSwitch_io_from_mat_0),
    .io_from_mat_1(ReadSwitch_io_from_mat_1),
    .io_from_mat_2(ReadSwitch_io_from_mat_2),
    .io_from_mat_3(ReadSwitch_io_from_mat_3),
    .io_from_mat_4(ReadSwitch_io_from_mat_4),
    .io_from_mat_5(ReadSwitch_io_from_mat_5),
    .io_from_mat_6(ReadSwitch_io_from_mat_6),
    .io_from_mat_7(ReadSwitch_io_from_mat_7),
    .io_from_mat_8(ReadSwitch_io_from_mat_8),
    .io_from_mat_9(ReadSwitch_io_from_mat_9),
    .io_from_mat_10(ReadSwitch_io_from_mat_10),
    .io_from_mat_11(ReadSwitch_io_from_mat_11),
    .io_from_mat_12(ReadSwitch_io_from_mat_12),
    .io_from_mat_13(ReadSwitch_io_from_mat_13),
    .io_from_mat_14(ReadSwitch_io_from_mat_14),
    .io_from_mat_15(ReadSwitch_io_from_mat_15),
    .io_from_mat_16(ReadSwitch_io_from_mat_16),
    .io_from_mat_17(ReadSwitch_io_from_mat_17),
    .io_from_mat_18(ReadSwitch_io_from_mat_18),
    .io_from_mat_19(ReadSwitch_io_from_mat_19),
    .io_from_mat_20(ReadSwitch_io_from_mat_20),
    .io_from_mat_21(ReadSwitch_io_from_mat_21),
    .io_from_mat_22(ReadSwitch_io_from_mat_22),
    .io_from_mat_23(ReadSwitch_io_from_mat_23),
    .io_from_mat_24(ReadSwitch_io_from_mat_24),
    .io_from_mat_25(ReadSwitch_io_from_mat_25),
    .io_from_mat_26(ReadSwitch_io_from_mat_26),
    .io_from_mat_27(ReadSwitch_io_from_mat_27),
    .io_from_mat_28(ReadSwitch_io_from_mat_28),
    .io_from_mat_29(ReadSwitch_io_from_mat_29),
    .io_from_mat_30(ReadSwitch_io_from_mat_30),
    .io_from_mat_31(ReadSwitch_io_from_mat_31),
    .io_from_mat_32(ReadSwitch_io_from_mat_32),
    .io_from_mat_33(ReadSwitch_io_from_mat_33),
    .io_from_mat_34(ReadSwitch_io_from_mat_34),
    .io_from_mat_35(ReadSwitch_io_from_mat_35),
    .io_from_mat_36(ReadSwitch_io_from_mat_36),
    .io_from_mat_37(ReadSwitch_io_from_mat_37),
    .io_from_mat_38(ReadSwitch_io_from_mat_38),
    .io_from_mat_39(ReadSwitch_io_from_mat_39),
    .io_from_mat_40(ReadSwitch_io_from_mat_40),
    .io_from_mat_41(ReadSwitch_io_from_mat_41),
    .io_from_mat_42(ReadSwitch_io_from_mat_42),
    .io_from_mat_43(ReadSwitch_io_from_mat_43),
    .io_from_mat_44(ReadSwitch_io_from_mat_44),
    .io_from_mat_45(ReadSwitch_io_from_mat_45),
    .io_from_mat_46(ReadSwitch_io_from_mat_46),
    .io_from_mat_47(ReadSwitch_io_from_mat_47),
    .io_from_mat_48(ReadSwitch_io_from_mat_48),
    .io_from_mat_49(ReadSwitch_io_from_mat_49),
    .io_from_mat_50(ReadSwitch_io_from_mat_50),
    .io_from_mat_51(ReadSwitch_io_from_mat_51),
    .io_from_mat_52(ReadSwitch_io_from_mat_52),
    .io_from_mat_53(ReadSwitch_io_from_mat_53),
    .io_from_mat_54(ReadSwitch_io_from_mat_54),
    .io_from_mat_55(ReadSwitch_io_from_mat_55),
    .io_from_mat_56(ReadSwitch_io_from_mat_56),
    .io_from_mat_57(ReadSwitch_io_from_mat_57),
    .io_from_mat_58(ReadSwitch_io_from_mat_58),
    .io_from_mat_59(ReadSwitch_io_from_mat_59),
    .io_from_mat_60(ReadSwitch_io_from_mat_60),
    .io_from_mat_61(ReadSwitch_io_from_mat_61),
    .io_from_mat_62(ReadSwitch_io_from_mat_62),
    .io_from_mat_63(ReadSwitch_io_from_mat_63),
    .io_from_up_0(ReadSwitch_io_from_up_0),
    .io_from_up_1(ReadSwitch_io_from_up_1),
    .io_from_up_2(ReadSwitch_io_from_up_2),
    .io_from_up_3(ReadSwitch_io_from_up_3),
    .io_from_up_4(ReadSwitch_io_from_up_4),
    .io_from_up_5(ReadSwitch_io_from_up_5),
    .io_from_up_6(ReadSwitch_io_from_up_6),
    .io_from_up_7(ReadSwitch_io_from_up_7),
    .io_from_up_8(ReadSwitch_io_from_up_8),
    .io_from_up_9(ReadSwitch_io_from_up_9),
    .io_from_down_0(ReadSwitch_io_from_down_0),
    .io_from_down_1(ReadSwitch_io_from_down_1),
    .io_from_down_2(ReadSwitch_io_from_down_2),
    .io_from_down_3(ReadSwitch_io_from_down_3),
    .io_from_down_4(ReadSwitch_io_from_down_4),
    .io_from_down_5(ReadSwitch_io_from_down_5),
    .io_from_down_6(ReadSwitch_io_from_down_6),
    .io_from_down_7(ReadSwitch_io_from_down_7),
    .io_from_down_8(ReadSwitch_io_from_down_8),
    .io_from_down_9(ReadSwitch_io_from_down_9),
    .io_from_left_0(ReadSwitch_io_from_left_0),
    .io_from_left_1(ReadSwitch_io_from_left_1),
    .io_from_left_2(ReadSwitch_io_from_left_2),
    .io_from_left_3(ReadSwitch_io_from_left_3),
    .io_from_left_4(ReadSwitch_io_from_left_4),
    .io_from_left_5(ReadSwitch_io_from_left_5),
    .io_from_left_6(ReadSwitch_io_from_left_6),
    .io_from_left_7(ReadSwitch_io_from_left_7),
    .io_from_right_0(ReadSwitch_io_from_right_0),
    .io_from_right_1(ReadSwitch_io_from_right_1),
    .io_from_right_2(ReadSwitch_io_from_right_2),
    .io_from_right_3(ReadSwitch_io_from_right_3),
    .io_from_right_4(ReadSwitch_io_from_right_4),
    .io_from_right_5(ReadSwitch_io_from_right_5),
    .io_from_right_6(ReadSwitch_io_from_right_6),
    .io_from_right_7(ReadSwitch_io_from_right_7),
    .io_from_weight_0(ReadSwitch_io_from_weight_0),
    .io_from_weight_1(ReadSwitch_io_from_weight_1),
    .io_from_weight_2(ReadSwitch_io_from_weight_2),
    .io_from_weight_3(ReadSwitch_io_from_weight_3),
    .io_from_weight_4(ReadSwitch_io_from_weight_4),
    .io_from_weight_5(ReadSwitch_io_from_weight_5),
    .io_from_weight_6(ReadSwitch_io_from_weight_6),
    .io_from_weight_7(ReadSwitch_io_from_weight_7),
    .io_from_weight_8(ReadSwitch_io_from_weight_8),
    .io_to_calc8x8_mat_0(ReadSwitch_io_to_calc8x8_mat_0),
    .io_to_calc8x8_mat_1(ReadSwitch_io_to_calc8x8_mat_1),
    .io_to_calc8x8_mat_2(ReadSwitch_io_to_calc8x8_mat_2),
    .io_to_calc8x8_mat_3(ReadSwitch_io_to_calc8x8_mat_3),
    .io_to_calc8x8_mat_4(ReadSwitch_io_to_calc8x8_mat_4),
    .io_to_calc8x8_mat_5(ReadSwitch_io_to_calc8x8_mat_5),
    .io_to_calc8x8_mat_6(ReadSwitch_io_to_calc8x8_mat_6),
    .io_to_calc8x8_mat_7(ReadSwitch_io_to_calc8x8_mat_7),
    .io_to_calc8x8_mat_8(ReadSwitch_io_to_calc8x8_mat_8),
    .io_to_calc8x8_mat_9(ReadSwitch_io_to_calc8x8_mat_9),
    .io_to_calc8x8_mat_10(ReadSwitch_io_to_calc8x8_mat_10),
    .io_to_calc8x8_mat_11(ReadSwitch_io_to_calc8x8_mat_11),
    .io_to_calc8x8_mat_12(ReadSwitch_io_to_calc8x8_mat_12),
    .io_to_calc8x8_mat_13(ReadSwitch_io_to_calc8x8_mat_13),
    .io_to_calc8x8_mat_14(ReadSwitch_io_to_calc8x8_mat_14),
    .io_to_calc8x8_mat_15(ReadSwitch_io_to_calc8x8_mat_15),
    .io_to_calc8x8_mat_16(ReadSwitch_io_to_calc8x8_mat_16),
    .io_to_calc8x8_mat_17(ReadSwitch_io_to_calc8x8_mat_17),
    .io_to_calc8x8_mat_18(ReadSwitch_io_to_calc8x8_mat_18),
    .io_to_calc8x8_mat_19(ReadSwitch_io_to_calc8x8_mat_19),
    .io_to_calc8x8_mat_20(ReadSwitch_io_to_calc8x8_mat_20),
    .io_to_calc8x8_mat_21(ReadSwitch_io_to_calc8x8_mat_21),
    .io_to_calc8x8_mat_22(ReadSwitch_io_to_calc8x8_mat_22),
    .io_to_calc8x8_mat_23(ReadSwitch_io_to_calc8x8_mat_23),
    .io_to_calc8x8_mat_24(ReadSwitch_io_to_calc8x8_mat_24),
    .io_to_calc8x8_mat_25(ReadSwitch_io_to_calc8x8_mat_25),
    .io_to_calc8x8_mat_26(ReadSwitch_io_to_calc8x8_mat_26),
    .io_to_calc8x8_mat_27(ReadSwitch_io_to_calc8x8_mat_27),
    .io_to_calc8x8_mat_28(ReadSwitch_io_to_calc8x8_mat_28),
    .io_to_calc8x8_mat_29(ReadSwitch_io_to_calc8x8_mat_29),
    .io_to_calc8x8_mat_30(ReadSwitch_io_to_calc8x8_mat_30),
    .io_to_calc8x8_mat_31(ReadSwitch_io_to_calc8x8_mat_31),
    .io_to_calc8x8_mat_32(ReadSwitch_io_to_calc8x8_mat_32),
    .io_to_calc8x8_mat_33(ReadSwitch_io_to_calc8x8_mat_33),
    .io_to_calc8x8_mat_34(ReadSwitch_io_to_calc8x8_mat_34),
    .io_to_calc8x8_mat_35(ReadSwitch_io_to_calc8x8_mat_35),
    .io_to_calc8x8_mat_36(ReadSwitch_io_to_calc8x8_mat_36),
    .io_to_calc8x8_mat_37(ReadSwitch_io_to_calc8x8_mat_37),
    .io_to_calc8x8_mat_38(ReadSwitch_io_to_calc8x8_mat_38),
    .io_to_calc8x8_mat_39(ReadSwitch_io_to_calc8x8_mat_39),
    .io_to_calc8x8_mat_40(ReadSwitch_io_to_calc8x8_mat_40),
    .io_to_calc8x8_mat_41(ReadSwitch_io_to_calc8x8_mat_41),
    .io_to_calc8x8_mat_42(ReadSwitch_io_to_calc8x8_mat_42),
    .io_to_calc8x8_mat_43(ReadSwitch_io_to_calc8x8_mat_43),
    .io_to_calc8x8_mat_44(ReadSwitch_io_to_calc8x8_mat_44),
    .io_to_calc8x8_mat_45(ReadSwitch_io_to_calc8x8_mat_45),
    .io_to_calc8x8_mat_46(ReadSwitch_io_to_calc8x8_mat_46),
    .io_to_calc8x8_mat_47(ReadSwitch_io_to_calc8x8_mat_47),
    .io_to_calc8x8_mat_48(ReadSwitch_io_to_calc8x8_mat_48),
    .io_to_calc8x8_mat_49(ReadSwitch_io_to_calc8x8_mat_49),
    .io_to_calc8x8_mat_50(ReadSwitch_io_to_calc8x8_mat_50),
    .io_to_calc8x8_mat_51(ReadSwitch_io_to_calc8x8_mat_51),
    .io_to_calc8x8_mat_52(ReadSwitch_io_to_calc8x8_mat_52),
    .io_to_calc8x8_mat_53(ReadSwitch_io_to_calc8x8_mat_53),
    .io_to_calc8x8_mat_54(ReadSwitch_io_to_calc8x8_mat_54),
    .io_to_calc8x8_mat_55(ReadSwitch_io_to_calc8x8_mat_55),
    .io_to_calc8x8_mat_56(ReadSwitch_io_to_calc8x8_mat_56),
    .io_to_calc8x8_mat_57(ReadSwitch_io_to_calc8x8_mat_57),
    .io_to_calc8x8_mat_58(ReadSwitch_io_to_calc8x8_mat_58),
    .io_to_calc8x8_mat_59(ReadSwitch_io_to_calc8x8_mat_59),
    .io_to_calc8x8_mat_60(ReadSwitch_io_to_calc8x8_mat_60),
    .io_to_calc8x8_mat_61(ReadSwitch_io_to_calc8x8_mat_61),
    .io_to_calc8x8_mat_62(ReadSwitch_io_to_calc8x8_mat_62),
    .io_to_calc8x8_mat_63(ReadSwitch_io_to_calc8x8_mat_63),
    .io_to_calc8x8_up_0(ReadSwitch_io_to_calc8x8_up_0),
    .io_to_calc8x8_up_1(ReadSwitch_io_to_calc8x8_up_1),
    .io_to_calc8x8_up_2(ReadSwitch_io_to_calc8x8_up_2),
    .io_to_calc8x8_up_3(ReadSwitch_io_to_calc8x8_up_3),
    .io_to_calc8x8_up_4(ReadSwitch_io_to_calc8x8_up_4),
    .io_to_calc8x8_up_5(ReadSwitch_io_to_calc8x8_up_5),
    .io_to_calc8x8_up_6(ReadSwitch_io_to_calc8x8_up_6),
    .io_to_calc8x8_up_7(ReadSwitch_io_to_calc8x8_up_7),
    .io_to_calc8x8_up_8(ReadSwitch_io_to_calc8x8_up_8),
    .io_to_calc8x8_up_9(ReadSwitch_io_to_calc8x8_up_9),
    .io_to_calc8x8_down_0(ReadSwitch_io_to_calc8x8_down_0),
    .io_to_calc8x8_down_1(ReadSwitch_io_to_calc8x8_down_1),
    .io_to_calc8x8_down_2(ReadSwitch_io_to_calc8x8_down_2),
    .io_to_calc8x8_down_3(ReadSwitch_io_to_calc8x8_down_3),
    .io_to_calc8x8_down_4(ReadSwitch_io_to_calc8x8_down_4),
    .io_to_calc8x8_down_5(ReadSwitch_io_to_calc8x8_down_5),
    .io_to_calc8x8_down_6(ReadSwitch_io_to_calc8x8_down_6),
    .io_to_calc8x8_down_7(ReadSwitch_io_to_calc8x8_down_7),
    .io_to_calc8x8_down_8(ReadSwitch_io_to_calc8x8_down_8),
    .io_to_calc8x8_down_9(ReadSwitch_io_to_calc8x8_down_9),
    .io_to_calc8x8_left_0(ReadSwitch_io_to_calc8x8_left_0),
    .io_to_calc8x8_left_1(ReadSwitch_io_to_calc8x8_left_1),
    .io_to_calc8x8_left_2(ReadSwitch_io_to_calc8x8_left_2),
    .io_to_calc8x8_left_3(ReadSwitch_io_to_calc8x8_left_3),
    .io_to_calc8x8_left_4(ReadSwitch_io_to_calc8x8_left_4),
    .io_to_calc8x8_left_5(ReadSwitch_io_to_calc8x8_left_5),
    .io_to_calc8x8_left_6(ReadSwitch_io_to_calc8x8_left_6),
    .io_to_calc8x8_left_7(ReadSwitch_io_to_calc8x8_left_7),
    .io_to_calc8x8_right_0(ReadSwitch_io_to_calc8x8_right_0),
    .io_to_calc8x8_right_1(ReadSwitch_io_to_calc8x8_right_1),
    .io_to_calc8x8_right_2(ReadSwitch_io_to_calc8x8_right_2),
    .io_to_calc8x8_right_3(ReadSwitch_io_to_calc8x8_right_3),
    .io_to_calc8x8_right_4(ReadSwitch_io_to_calc8x8_right_4),
    .io_to_calc8x8_right_5(ReadSwitch_io_to_calc8x8_right_5),
    .io_to_calc8x8_right_6(ReadSwitch_io_to_calc8x8_right_6),
    .io_to_calc8x8_right_7(ReadSwitch_io_to_calc8x8_right_7),
    .io_to_weight_0_real_0(ReadSwitch_io_to_weight_0_real_0),
    .io_to_weight_0_real_1(ReadSwitch_io_to_weight_0_real_1),
    .io_to_weight_0_real_2(ReadSwitch_io_to_weight_0_real_2),
    .io_to_weight_0_real_3(ReadSwitch_io_to_weight_0_real_3),
    .io_to_weight_0_real_4(ReadSwitch_io_to_weight_0_real_4),
    .io_to_weight_0_real_5(ReadSwitch_io_to_weight_0_real_5),
    .io_to_weight_0_real_6(ReadSwitch_io_to_weight_0_real_6),
    .io_to_weight_0_real_7(ReadSwitch_io_to_weight_0_real_7),
    .io_to_weight_0_real_8(ReadSwitch_io_to_weight_0_real_8),
    .io_to_weight_0_real_9(ReadSwitch_io_to_weight_0_real_9),
    .io_to_weight_0_real_10(ReadSwitch_io_to_weight_0_real_10),
    .io_to_weight_0_real_11(ReadSwitch_io_to_weight_0_real_11),
    .io_to_weight_0_real_12(ReadSwitch_io_to_weight_0_real_12),
    .io_to_weight_0_real_13(ReadSwitch_io_to_weight_0_real_13),
    .io_to_weight_0_real_14(ReadSwitch_io_to_weight_0_real_14),
    .io_to_weight_0_real_15(ReadSwitch_io_to_weight_0_real_15),
    .io_to_weight_1_real_0(ReadSwitch_io_to_weight_1_real_0),
    .io_to_weight_1_real_1(ReadSwitch_io_to_weight_1_real_1),
    .io_to_weight_1_real_2(ReadSwitch_io_to_weight_1_real_2),
    .io_to_weight_1_real_3(ReadSwitch_io_to_weight_1_real_3),
    .io_to_weight_1_real_4(ReadSwitch_io_to_weight_1_real_4),
    .io_to_weight_1_real_5(ReadSwitch_io_to_weight_1_real_5),
    .io_to_weight_1_real_6(ReadSwitch_io_to_weight_1_real_6),
    .io_to_weight_1_real_7(ReadSwitch_io_to_weight_1_real_7),
    .io_to_weight_1_real_8(ReadSwitch_io_to_weight_1_real_8),
    .io_to_weight_1_real_9(ReadSwitch_io_to_weight_1_real_9),
    .io_to_weight_1_real_10(ReadSwitch_io_to_weight_1_real_10),
    .io_to_weight_1_real_11(ReadSwitch_io_to_weight_1_real_11),
    .io_to_weight_1_real_12(ReadSwitch_io_to_weight_1_real_12),
    .io_to_weight_1_real_13(ReadSwitch_io_to_weight_1_real_13),
    .io_to_weight_1_real_14(ReadSwitch_io_to_weight_1_real_14),
    .io_to_weight_1_real_15(ReadSwitch_io_to_weight_1_real_15),
    .io_to_weight_2_real_0(ReadSwitch_io_to_weight_2_real_0),
    .io_to_weight_2_real_1(ReadSwitch_io_to_weight_2_real_1),
    .io_to_weight_2_real_2(ReadSwitch_io_to_weight_2_real_2),
    .io_to_weight_2_real_3(ReadSwitch_io_to_weight_2_real_3),
    .io_to_weight_2_real_4(ReadSwitch_io_to_weight_2_real_4),
    .io_to_weight_2_real_5(ReadSwitch_io_to_weight_2_real_5),
    .io_to_weight_2_real_6(ReadSwitch_io_to_weight_2_real_6),
    .io_to_weight_2_real_7(ReadSwitch_io_to_weight_2_real_7),
    .io_to_weight_2_real_8(ReadSwitch_io_to_weight_2_real_8),
    .io_to_weight_2_real_9(ReadSwitch_io_to_weight_2_real_9),
    .io_to_weight_2_real_10(ReadSwitch_io_to_weight_2_real_10),
    .io_to_weight_2_real_11(ReadSwitch_io_to_weight_2_real_11),
    .io_to_weight_2_real_12(ReadSwitch_io_to_weight_2_real_12),
    .io_to_weight_2_real_13(ReadSwitch_io_to_weight_2_real_13),
    .io_to_weight_2_real_14(ReadSwitch_io_to_weight_2_real_14),
    .io_to_weight_2_real_15(ReadSwitch_io_to_weight_2_real_15),
    .io_to_weight_3_real_0(ReadSwitch_io_to_weight_3_real_0),
    .io_to_weight_3_real_1(ReadSwitch_io_to_weight_3_real_1),
    .io_to_weight_3_real_2(ReadSwitch_io_to_weight_3_real_2),
    .io_to_weight_3_real_3(ReadSwitch_io_to_weight_3_real_3),
    .io_to_weight_3_real_4(ReadSwitch_io_to_weight_3_real_4),
    .io_to_weight_3_real_5(ReadSwitch_io_to_weight_3_real_5),
    .io_to_weight_3_real_6(ReadSwitch_io_to_weight_3_real_6),
    .io_to_weight_3_real_7(ReadSwitch_io_to_weight_3_real_7),
    .io_to_weight_3_real_8(ReadSwitch_io_to_weight_3_real_8),
    .io_to_weight_3_real_9(ReadSwitch_io_to_weight_3_real_9),
    .io_to_weight_3_real_10(ReadSwitch_io_to_weight_3_real_10),
    .io_to_weight_3_real_11(ReadSwitch_io_to_weight_3_real_11),
    .io_to_weight_3_real_12(ReadSwitch_io_to_weight_3_real_12),
    .io_to_weight_3_real_13(ReadSwitch_io_to_weight_3_real_13),
    .io_to_weight_3_real_14(ReadSwitch_io_to_weight_3_real_14),
    .io_to_weight_3_real_15(ReadSwitch_io_to_weight_3_real_15)
  );
  WeightReader WeightReader ( // @[top.scala 18:29]
    .clock(WeightReader_clock),
    .reset(WeightReader_reset),
    .io_valid_in(WeightReader_io_valid_in),
    .io_flag_job(WeightReader_io_flag_job),
    .io_addr_end(WeightReader_io_addr_end),
    .io_addr(WeightReader_io_addr)
  );
  Calc8x8 Calc8x8 ( // @[top.scala 19:25]
    .clock(Calc8x8_clock),
    .reset(Calc8x8_reset),
    .io_input_mat_0(Calc8x8_io_input_mat_0),
    .io_input_mat_1(Calc8x8_io_input_mat_1),
    .io_input_mat_2(Calc8x8_io_input_mat_2),
    .io_input_mat_3(Calc8x8_io_input_mat_3),
    .io_input_mat_4(Calc8x8_io_input_mat_4),
    .io_input_mat_5(Calc8x8_io_input_mat_5),
    .io_input_mat_6(Calc8x8_io_input_mat_6),
    .io_input_mat_7(Calc8x8_io_input_mat_7),
    .io_input_mat_8(Calc8x8_io_input_mat_8),
    .io_input_mat_9(Calc8x8_io_input_mat_9),
    .io_input_mat_10(Calc8x8_io_input_mat_10),
    .io_input_mat_11(Calc8x8_io_input_mat_11),
    .io_input_mat_12(Calc8x8_io_input_mat_12),
    .io_input_mat_13(Calc8x8_io_input_mat_13),
    .io_input_mat_14(Calc8x8_io_input_mat_14),
    .io_input_mat_15(Calc8x8_io_input_mat_15),
    .io_input_mat_16(Calc8x8_io_input_mat_16),
    .io_input_mat_17(Calc8x8_io_input_mat_17),
    .io_input_mat_18(Calc8x8_io_input_mat_18),
    .io_input_mat_19(Calc8x8_io_input_mat_19),
    .io_input_mat_20(Calc8x8_io_input_mat_20),
    .io_input_mat_21(Calc8x8_io_input_mat_21),
    .io_input_mat_22(Calc8x8_io_input_mat_22),
    .io_input_mat_23(Calc8x8_io_input_mat_23),
    .io_input_mat_24(Calc8x8_io_input_mat_24),
    .io_input_mat_25(Calc8x8_io_input_mat_25),
    .io_input_mat_26(Calc8x8_io_input_mat_26),
    .io_input_mat_27(Calc8x8_io_input_mat_27),
    .io_input_mat_28(Calc8x8_io_input_mat_28),
    .io_input_mat_29(Calc8x8_io_input_mat_29),
    .io_input_mat_30(Calc8x8_io_input_mat_30),
    .io_input_mat_31(Calc8x8_io_input_mat_31),
    .io_input_mat_32(Calc8x8_io_input_mat_32),
    .io_input_mat_33(Calc8x8_io_input_mat_33),
    .io_input_mat_34(Calc8x8_io_input_mat_34),
    .io_input_mat_35(Calc8x8_io_input_mat_35),
    .io_input_mat_36(Calc8x8_io_input_mat_36),
    .io_input_mat_37(Calc8x8_io_input_mat_37),
    .io_input_mat_38(Calc8x8_io_input_mat_38),
    .io_input_mat_39(Calc8x8_io_input_mat_39),
    .io_input_mat_40(Calc8x8_io_input_mat_40),
    .io_input_mat_41(Calc8x8_io_input_mat_41),
    .io_input_mat_42(Calc8x8_io_input_mat_42),
    .io_input_mat_43(Calc8x8_io_input_mat_43),
    .io_input_mat_44(Calc8x8_io_input_mat_44),
    .io_input_mat_45(Calc8x8_io_input_mat_45),
    .io_input_mat_46(Calc8x8_io_input_mat_46),
    .io_input_mat_47(Calc8x8_io_input_mat_47),
    .io_input_mat_48(Calc8x8_io_input_mat_48),
    .io_input_mat_49(Calc8x8_io_input_mat_49),
    .io_input_mat_50(Calc8x8_io_input_mat_50),
    .io_input_mat_51(Calc8x8_io_input_mat_51),
    .io_input_mat_52(Calc8x8_io_input_mat_52),
    .io_input_mat_53(Calc8x8_io_input_mat_53),
    .io_input_mat_54(Calc8x8_io_input_mat_54),
    .io_input_mat_55(Calc8x8_io_input_mat_55),
    .io_input_mat_56(Calc8x8_io_input_mat_56),
    .io_input_mat_57(Calc8x8_io_input_mat_57),
    .io_input_mat_58(Calc8x8_io_input_mat_58),
    .io_input_mat_59(Calc8x8_io_input_mat_59),
    .io_input_mat_60(Calc8x8_io_input_mat_60),
    .io_input_mat_61(Calc8x8_io_input_mat_61),
    .io_input_mat_62(Calc8x8_io_input_mat_62),
    .io_input_mat_63(Calc8x8_io_input_mat_63),
    .io_input_up_0(Calc8x8_io_input_up_0),
    .io_input_up_1(Calc8x8_io_input_up_1),
    .io_input_up_2(Calc8x8_io_input_up_2),
    .io_input_up_3(Calc8x8_io_input_up_3),
    .io_input_up_4(Calc8x8_io_input_up_4),
    .io_input_up_5(Calc8x8_io_input_up_5),
    .io_input_up_6(Calc8x8_io_input_up_6),
    .io_input_up_7(Calc8x8_io_input_up_7),
    .io_input_up_8(Calc8x8_io_input_up_8),
    .io_input_up_9(Calc8x8_io_input_up_9),
    .io_input_down_0(Calc8x8_io_input_down_0),
    .io_input_down_1(Calc8x8_io_input_down_1),
    .io_input_down_2(Calc8x8_io_input_down_2),
    .io_input_down_3(Calc8x8_io_input_down_3),
    .io_input_down_4(Calc8x8_io_input_down_4),
    .io_input_down_5(Calc8x8_io_input_down_5),
    .io_input_down_6(Calc8x8_io_input_down_6),
    .io_input_down_7(Calc8x8_io_input_down_7),
    .io_input_down_8(Calc8x8_io_input_down_8),
    .io_input_down_9(Calc8x8_io_input_down_9),
    .io_input_left_0(Calc8x8_io_input_left_0),
    .io_input_left_1(Calc8x8_io_input_left_1),
    .io_input_left_2(Calc8x8_io_input_left_2),
    .io_input_left_3(Calc8x8_io_input_left_3),
    .io_input_left_4(Calc8x8_io_input_left_4),
    .io_input_left_5(Calc8x8_io_input_left_5),
    .io_input_left_6(Calc8x8_io_input_left_6),
    .io_input_left_7(Calc8x8_io_input_left_7),
    .io_input_right_0(Calc8x8_io_input_right_0),
    .io_input_right_1(Calc8x8_io_input_right_1),
    .io_input_right_2(Calc8x8_io_input_right_2),
    .io_input_right_3(Calc8x8_io_input_right_3),
    .io_input_right_4(Calc8x8_io_input_right_4),
    .io_input_right_5(Calc8x8_io_input_right_5),
    .io_input_right_6(Calc8x8_io_input_right_6),
    .io_input_right_7(Calc8x8_io_input_right_7),
    .io_flag(Calc8x8_io_flag),
    .io_weight_0_real_0(Calc8x8_io_weight_0_real_0),
    .io_weight_0_real_1(Calc8x8_io_weight_0_real_1),
    .io_weight_0_real_2(Calc8x8_io_weight_0_real_2),
    .io_weight_0_real_3(Calc8x8_io_weight_0_real_3),
    .io_weight_0_real_4(Calc8x8_io_weight_0_real_4),
    .io_weight_0_real_5(Calc8x8_io_weight_0_real_5),
    .io_weight_0_real_6(Calc8x8_io_weight_0_real_6),
    .io_weight_0_real_7(Calc8x8_io_weight_0_real_7),
    .io_weight_0_real_8(Calc8x8_io_weight_0_real_8),
    .io_weight_0_real_9(Calc8x8_io_weight_0_real_9),
    .io_weight_0_real_10(Calc8x8_io_weight_0_real_10),
    .io_weight_0_real_11(Calc8x8_io_weight_0_real_11),
    .io_weight_0_real_12(Calc8x8_io_weight_0_real_12),
    .io_weight_0_real_13(Calc8x8_io_weight_0_real_13),
    .io_weight_0_real_14(Calc8x8_io_weight_0_real_14),
    .io_weight_0_real_15(Calc8x8_io_weight_0_real_15),
    .io_weight_1_real_0(Calc8x8_io_weight_1_real_0),
    .io_weight_1_real_1(Calc8x8_io_weight_1_real_1),
    .io_weight_1_real_2(Calc8x8_io_weight_1_real_2),
    .io_weight_1_real_3(Calc8x8_io_weight_1_real_3),
    .io_weight_1_real_4(Calc8x8_io_weight_1_real_4),
    .io_weight_1_real_5(Calc8x8_io_weight_1_real_5),
    .io_weight_1_real_6(Calc8x8_io_weight_1_real_6),
    .io_weight_1_real_7(Calc8x8_io_weight_1_real_7),
    .io_weight_1_real_8(Calc8x8_io_weight_1_real_8),
    .io_weight_1_real_9(Calc8x8_io_weight_1_real_9),
    .io_weight_1_real_10(Calc8x8_io_weight_1_real_10),
    .io_weight_1_real_11(Calc8x8_io_weight_1_real_11),
    .io_weight_1_real_12(Calc8x8_io_weight_1_real_12),
    .io_weight_1_real_13(Calc8x8_io_weight_1_real_13),
    .io_weight_1_real_14(Calc8x8_io_weight_1_real_14),
    .io_weight_1_real_15(Calc8x8_io_weight_1_real_15),
    .io_weight_2_real_0(Calc8x8_io_weight_2_real_0),
    .io_weight_2_real_1(Calc8x8_io_weight_2_real_1),
    .io_weight_2_real_2(Calc8x8_io_weight_2_real_2),
    .io_weight_2_real_3(Calc8x8_io_weight_2_real_3),
    .io_weight_2_real_4(Calc8x8_io_weight_2_real_4),
    .io_weight_2_real_5(Calc8x8_io_weight_2_real_5),
    .io_weight_2_real_6(Calc8x8_io_weight_2_real_6),
    .io_weight_2_real_7(Calc8x8_io_weight_2_real_7),
    .io_weight_2_real_8(Calc8x8_io_weight_2_real_8),
    .io_weight_2_real_9(Calc8x8_io_weight_2_real_9),
    .io_weight_2_real_10(Calc8x8_io_weight_2_real_10),
    .io_weight_2_real_11(Calc8x8_io_weight_2_real_11),
    .io_weight_2_real_12(Calc8x8_io_weight_2_real_12),
    .io_weight_2_real_13(Calc8x8_io_weight_2_real_13),
    .io_weight_2_real_14(Calc8x8_io_weight_2_real_14),
    .io_weight_2_real_15(Calc8x8_io_weight_2_real_15),
    .io_weight_3_real_0(Calc8x8_io_weight_3_real_0),
    .io_weight_3_real_1(Calc8x8_io_weight_3_real_1),
    .io_weight_3_real_2(Calc8x8_io_weight_3_real_2),
    .io_weight_3_real_3(Calc8x8_io_weight_3_real_3),
    .io_weight_3_real_4(Calc8x8_io_weight_3_real_4),
    .io_weight_3_real_5(Calc8x8_io_weight_3_real_5),
    .io_weight_3_real_6(Calc8x8_io_weight_3_real_6),
    .io_weight_3_real_7(Calc8x8_io_weight_3_real_7),
    .io_weight_3_real_8(Calc8x8_io_weight_3_real_8),
    .io_weight_3_real_9(Calc8x8_io_weight_3_real_9),
    .io_weight_3_real_10(Calc8x8_io_weight_3_real_10),
    .io_weight_3_real_11(Calc8x8_io_weight_3_real_11),
    .io_weight_3_real_12(Calc8x8_io_weight_3_real_12),
    .io_weight_3_real_13(Calc8x8_io_weight_3_real_13),
    .io_weight_3_real_14(Calc8x8_io_weight_3_real_14),
    .io_weight_3_real_15(Calc8x8_io_weight_3_real_15),
    .io_output_mat_0(Calc8x8_io_output_mat_0),
    .io_output_mat_1(Calc8x8_io_output_mat_1),
    .io_output_mat_2(Calc8x8_io_output_mat_2),
    .io_output_mat_3(Calc8x8_io_output_mat_3),
    .io_output_mat_4(Calc8x8_io_output_mat_4),
    .io_output_mat_5(Calc8x8_io_output_mat_5),
    .io_output_mat_6(Calc8x8_io_output_mat_6),
    .io_output_mat_7(Calc8x8_io_output_mat_7),
    .io_output_mat_8(Calc8x8_io_output_mat_8),
    .io_output_mat_9(Calc8x8_io_output_mat_9),
    .io_output_mat_10(Calc8x8_io_output_mat_10),
    .io_output_mat_11(Calc8x8_io_output_mat_11),
    .io_output_mat_12(Calc8x8_io_output_mat_12),
    .io_output_mat_13(Calc8x8_io_output_mat_13),
    .io_output_mat_14(Calc8x8_io_output_mat_14),
    .io_output_mat_15(Calc8x8_io_output_mat_15),
    .io_output_mat_16(Calc8x8_io_output_mat_16),
    .io_output_mat_17(Calc8x8_io_output_mat_17),
    .io_output_mat_18(Calc8x8_io_output_mat_18),
    .io_output_mat_19(Calc8x8_io_output_mat_19),
    .io_output_mat_20(Calc8x8_io_output_mat_20),
    .io_output_mat_21(Calc8x8_io_output_mat_21),
    .io_output_mat_22(Calc8x8_io_output_mat_22),
    .io_output_mat_23(Calc8x8_io_output_mat_23),
    .io_output_mat_24(Calc8x8_io_output_mat_24),
    .io_output_mat_25(Calc8x8_io_output_mat_25),
    .io_output_mat_26(Calc8x8_io_output_mat_26),
    .io_output_mat_27(Calc8x8_io_output_mat_27),
    .io_output_mat_28(Calc8x8_io_output_mat_28),
    .io_output_mat_29(Calc8x8_io_output_mat_29),
    .io_output_mat_30(Calc8x8_io_output_mat_30),
    .io_output_mat_31(Calc8x8_io_output_mat_31),
    .io_output_mat_32(Calc8x8_io_output_mat_32),
    .io_output_mat_33(Calc8x8_io_output_mat_33),
    .io_output_mat_34(Calc8x8_io_output_mat_34),
    .io_output_mat_35(Calc8x8_io_output_mat_35),
    .io_output_mat_36(Calc8x8_io_output_mat_36),
    .io_output_mat_37(Calc8x8_io_output_mat_37),
    .io_output_mat_38(Calc8x8_io_output_mat_38),
    .io_output_mat_39(Calc8x8_io_output_mat_39),
    .io_output_mat_40(Calc8x8_io_output_mat_40),
    .io_output_mat_41(Calc8x8_io_output_mat_41),
    .io_output_mat_42(Calc8x8_io_output_mat_42),
    .io_output_mat_43(Calc8x8_io_output_mat_43),
    .io_output_mat_44(Calc8x8_io_output_mat_44),
    .io_output_mat_45(Calc8x8_io_output_mat_45),
    .io_output_mat_46(Calc8x8_io_output_mat_46),
    .io_output_mat_47(Calc8x8_io_output_mat_47),
    .io_output_mat_48(Calc8x8_io_output_mat_48),
    .io_output_mat_49(Calc8x8_io_output_mat_49),
    .io_output_mat_50(Calc8x8_io_output_mat_50),
    .io_output_mat_51(Calc8x8_io_output_mat_51),
    .io_output_mat_52(Calc8x8_io_output_mat_52),
    .io_output_mat_53(Calc8x8_io_output_mat_53),
    .io_output_mat_54(Calc8x8_io_output_mat_54),
    .io_output_mat_55(Calc8x8_io_output_mat_55),
    .io_output_mat_56(Calc8x8_io_output_mat_56),
    .io_output_mat_57(Calc8x8_io_output_mat_57),
    .io_output_mat_58(Calc8x8_io_output_mat_58),
    .io_output_mat_59(Calc8x8_io_output_mat_59),
    .io_output_mat_60(Calc8x8_io_output_mat_60),
    .io_output_mat_61(Calc8x8_io_output_mat_61),
    .io_output_mat_62(Calc8x8_io_output_mat_62),
    .io_output_mat_63(Calc8x8_io_output_mat_63),
    .io_valid_in(Calc8x8_io_valid_in),
    .io_valid_out(Calc8x8_io_valid_out)
  );
  Accumu Accumu ( // @[top.scala 20:22]
    .clock(Accumu_clock),
    .reset(Accumu_reset),
    .io_valid_in(Accumu_io_valid_in),
    .io_valid_out(Accumu_io_valid_out),
    .io_flag_job(Accumu_io_flag_job),
    .io_in_from_calc8x8_mat_0(Accumu_io_in_from_calc8x8_mat_0),
    .io_in_from_calc8x8_mat_1(Accumu_io_in_from_calc8x8_mat_1),
    .io_in_from_calc8x8_mat_2(Accumu_io_in_from_calc8x8_mat_2),
    .io_in_from_calc8x8_mat_3(Accumu_io_in_from_calc8x8_mat_3),
    .io_in_from_calc8x8_mat_4(Accumu_io_in_from_calc8x8_mat_4),
    .io_in_from_calc8x8_mat_5(Accumu_io_in_from_calc8x8_mat_5),
    .io_in_from_calc8x8_mat_6(Accumu_io_in_from_calc8x8_mat_6),
    .io_in_from_calc8x8_mat_7(Accumu_io_in_from_calc8x8_mat_7),
    .io_in_from_calc8x8_mat_8(Accumu_io_in_from_calc8x8_mat_8),
    .io_in_from_calc8x8_mat_9(Accumu_io_in_from_calc8x8_mat_9),
    .io_in_from_calc8x8_mat_10(Accumu_io_in_from_calc8x8_mat_10),
    .io_in_from_calc8x8_mat_11(Accumu_io_in_from_calc8x8_mat_11),
    .io_in_from_calc8x8_mat_12(Accumu_io_in_from_calc8x8_mat_12),
    .io_in_from_calc8x8_mat_13(Accumu_io_in_from_calc8x8_mat_13),
    .io_in_from_calc8x8_mat_14(Accumu_io_in_from_calc8x8_mat_14),
    .io_in_from_calc8x8_mat_15(Accumu_io_in_from_calc8x8_mat_15),
    .io_in_from_calc8x8_mat_16(Accumu_io_in_from_calc8x8_mat_16),
    .io_in_from_calc8x8_mat_17(Accumu_io_in_from_calc8x8_mat_17),
    .io_in_from_calc8x8_mat_18(Accumu_io_in_from_calc8x8_mat_18),
    .io_in_from_calc8x8_mat_19(Accumu_io_in_from_calc8x8_mat_19),
    .io_in_from_calc8x8_mat_20(Accumu_io_in_from_calc8x8_mat_20),
    .io_in_from_calc8x8_mat_21(Accumu_io_in_from_calc8x8_mat_21),
    .io_in_from_calc8x8_mat_22(Accumu_io_in_from_calc8x8_mat_22),
    .io_in_from_calc8x8_mat_23(Accumu_io_in_from_calc8x8_mat_23),
    .io_in_from_calc8x8_mat_24(Accumu_io_in_from_calc8x8_mat_24),
    .io_in_from_calc8x8_mat_25(Accumu_io_in_from_calc8x8_mat_25),
    .io_in_from_calc8x8_mat_26(Accumu_io_in_from_calc8x8_mat_26),
    .io_in_from_calc8x8_mat_27(Accumu_io_in_from_calc8x8_mat_27),
    .io_in_from_calc8x8_mat_28(Accumu_io_in_from_calc8x8_mat_28),
    .io_in_from_calc8x8_mat_29(Accumu_io_in_from_calc8x8_mat_29),
    .io_in_from_calc8x8_mat_30(Accumu_io_in_from_calc8x8_mat_30),
    .io_in_from_calc8x8_mat_31(Accumu_io_in_from_calc8x8_mat_31),
    .io_in_from_calc8x8_mat_32(Accumu_io_in_from_calc8x8_mat_32),
    .io_in_from_calc8x8_mat_33(Accumu_io_in_from_calc8x8_mat_33),
    .io_in_from_calc8x8_mat_34(Accumu_io_in_from_calc8x8_mat_34),
    .io_in_from_calc8x8_mat_35(Accumu_io_in_from_calc8x8_mat_35),
    .io_in_from_calc8x8_mat_36(Accumu_io_in_from_calc8x8_mat_36),
    .io_in_from_calc8x8_mat_37(Accumu_io_in_from_calc8x8_mat_37),
    .io_in_from_calc8x8_mat_38(Accumu_io_in_from_calc8x8_mat_38),
    .io_in_from_calc8x8_mat_39(Accumu_io_in_from_calc8x8_mat_39),
    .io_in_from_calc8x8_mat_40(Accumu_io_in_from_calc8x8_mat_40),
    .io_in_from_calc8x8_mat_41(Accumu_io_in_from_calc8x8_mat_41),
    .io_in_from_calc8x8_mat_42(Accumu_io_in_from_calc8x8_mat_42),
    .io_in_from_calc8x8_mat_43(Accumu_io_in_from_calc8x8_mat_43),
    .io_in_from_calc8x8_mat_44(Accumu_io_in_from_calc8x8_mat_44),
    .io_in_from_calc8x8_mat_45(Accumu_io_in_from_calc8x8_mat_45),
    .io_in_from_calc8x8_mat_46(Accumu_io_in_from_calc8x8_mat_46),
    .io_in_from_calc8x8_mat_47(Accumu_io_in_from_calc8x8_mat_47),
    .io_in_from_calc8x8_mat_48(Accumu_io_in_from_calc8x8_mat_48),
    .io_in_from_calc8x8_mat_49(Accumu_io_in_from_calc8x8_mat_49),
    .io_in_from_calc8x8_mat_50(Accumu_io_in_from_calc8x8_mat_50),
    .io_in_from_calc8x8_mat_51(Accumu_io_in_from_calc8x8_mat_51),
    .io_in_from_calc8x8_mat_52(Accumu_io_in_from_calc8x8_mat_52),
    .io_in_from_calc8x8_mat_53(Accumu_io_in_from_calc8x8_mat_53),
    .io_in_from_calc8x8_mat_54(Accumu_io_in_from_calc8x8_mat_54),
    .io_in_from_calc8x8_mat_55(Accumu_io_in_from_calc8x8_mat_55),
    .io_in_from_calc8x8_mat_56(Accumu_io_in_from_calc8x8_mat_56),
    .io_in_from_calc8x8_mat_57(Accumu_io_in_from_calc8x8_mat_57),
    .io_in_from_calc8x8_mat_58(Accumu_io_in_from_calc8x8_mat_58),
    .io_in_from_calc8x8_mat_59(Accumu_io_in_from_calc8x8_mat_59),
    .io_in_from_calc8x8_mat_60(Accumu_io_in_from_calc8x8_mat_60),
    .io_in_from_calc8x8_mat_61(Accumu_io_in_from_calc8x8_mat_61),
    .io_in_from_calc8x8_mat_62(Accumu_io_in_from_calc8x8_mat_62),
    .io_in_from_calc8x8_mat_63(Accumu_io_in_from_calc8x8_mat_63),
    .io_result_mat_0(Accumu_io_result_mat_0),
    .io_result_mat_1(Accumu_io_result_mat_1),
    .io_result_mat_2(Accumu_io_result_mat_2),
    .io_result_mat_3(Accumu_io_result_mat_3),
    .io_result_mat_4(Accumu_io_result_mat_4),
    .io_result_mat_5(Accumu_io_result_mat_5),
    .io_result_mat_6(Accumu_io_result_mat_6),
    .io_result_mat_7(Accumu_io_result_mat_7),
    .io_result_mat_8(Accumu_io_result_mat_8),
    .io_result_mat_9(Accumu_io_result_mat_9),
    .io_result_mat_10(Accumu_io_result_mat_10),
    .io_result_mat_11(Accumu_io_result_mat_11),
    .io_result_mat_12(Accumu_io_result_mat_12),
    .io_result_mat_13(Accumu_io_result_mat_13),
    .io_result_mat_14(Accumu_io_result_mat_14),
    .io_result_mat_15(Accumu_io_result_mat_15),
    .io_result_mat_16(Accumu_io_result_mat_16),
    .io_result_mat_17(Accumu_io_result_mat_17),
    .io_result_mat_18(Accumu_io_result_mat_18),
    .io_result_mat_19(Accumu_io_result_mat_19),
    .io_result_mat_20(Accumu_io_result_mat_20),
    .io_result_mat_21(Accumu_io_result_mat_21),
    .io_result_mat_22(Accumu_io_result_mat_22),
    .io_result_mat_23(Accumu_io_result_mat_23),
    .io_result_mat_24(Accumu_io_result_mat_24),
    .io_result_mat_25(Accumu_io_result_mat_25),
    .io_result_mat_26(Accumu_io_result_mat_26),
    .io_result_mat_27(Accumu_io_result_mat_27),
    .io_result_mat_28(Accumu_io_result_mat_28),
    .io_result_mat_29(Accumu_io_result_mat_29),
    .io_result_mat_30(Accumu_io_result_mat_30),
    .io_result_mat_31(Accumu_io_result_mat_31),
    .io_result_mat_32(Accumu_io_result_mat_32),
    .io_result_mat_33(Accumu_io_result_mat_33),
    .io_result_mat_34(Accumu_io_result_mat_34),
    .io_result_mat_35(Accumu_io_result_mat_35),
    .io_result_mat_36(Accumu_io_result_mat_36),
    .io_result_mat_37(Accumu_io_result_mat_37),
    .io_result_mat_38(Accumu_io_result_mat_38),
    .io_result_mat_39(Accumu_io_result_mat_39),
    .io_result_mat_40(Accumu_io_result_mat_40),
    .io_result_mat_41(Accumu_io_result_mat_41),
    .io_result_mat_42(Accumu_io_result_mat_42),
    .io_result_mat_43(Accumu_io_result_mat_43),
    .io_result_mat_44(Accumu_io_result_mat_44),
    .io_result_mat_45(Accumu_io_result_mat_45),
    .io_result_mat_46(Accumu_io_result_mat_46),
    .io_result_mat_47(Accumu_io_result_mat_47),
    .io_result_mat_48(Accumu_io_result_mat_48),
    .io_result_mat_49(Accumu_io_result_mat_49),
    .io_result_mat_50(Accumu_io_result_mat_50),
    .io_result_mat_51(Accumu_io_result_mat_51),
    .io_result_mat_52(Accumu_io_result_mat_52),
    .io_result_mat_53(Accumu_io_result_mat_53),
    .io_result_mat_54(Accumu_io_result_mat_54),
    .io_result_mat_55(Accumu_io_result_mat_55),
    .io_result_mat_56(Accumu_io_result_mat_56),
    .io_result_mat_57(Accumu_io_result_mat_57),
    .io_result_mat_58(Accumu_io_result_mat_58),
    .io_result_mat_59(Accumu_io_result_mat_59),
    .io_result_mat_60(Accumu_io_result_mat_60),
    .io_result_mat_61(Accumu_io_result_mat_61),
    .io_result_mat_62(Accumu_io_result_mat_62),
    .io_result_mat_63(Accumu_io_result_mat_63),
    .io_csum(Accumu_io_csum),
    .io_bias_end_addr(Accumu_io_bias_end_addr),
    .io_bias_addr(Accumu_io_bias_addr),
    .io_bias_in(Accumu_io_bias_in),
    .io_is_in_use(Accumu_io_is_in_use)
  );
  Quant Quant ( // @[top.scala 21:23]
    .clock(Quant_clock),
    .reset(Quant_reset),
    .io_valid_in(Quant_io_valid_in),
    .io_valid_out(Quant_io_valid_out),
    .io_flag_job(Quant_io_flag_job),
    .io_in_from_accumu_mat_0(Quant_io_in_from_accumu_mat_0),
    .io_in_from_accumu_mat_1(Quant_io_in_from_accumu_mat_1),
    .io_in_from_accumu_mat_2(Quant_io_in_from_accumu_mat_2),
    .io_in_from_accumu_mat_3(Quant_io_in_from_accumu_mat_3),
    .io_in_from_accumu_mat_4(Quant_io_in_from_accumu_mat_4),
    .io_in_from_accumu_mat_5(Quant_io_in_from_accumu_mat_5),
    .io_in_from_accumu_mat_6(Quant_io_in_from_accumu_mat_6),
    .io_in_from_accumu_mat_7(Quant_io_in_from_accumu_mat_7),
    .io_in_from_accumu_mat_8(Quant_io_in_from_accumu_mat_8),
    .io_in_from_accumu_mat_9(Quant_io_in_from_accumu_mat_9),
    .io_in_from_accumu_mat_10(Quant_io_in_from_accumu_mat_10),
    .io_in_from_accumu_mat_11(Quant_io_in_from_accumu_mat_11),
    .io_in_from_accumu_mat_12(Quant_io_in_from_accumu_mat_12),
    .io_in_from_accumu_mat_13(Quant_io_in_from_accumu_mat_13),
    .io_in_from_accumu_mat_14(Quant_io_in_from_accumu_mat_14),
    .io_in_from_accumu_mat_15(Quant_io_in_from_accumu_mat_15),
    .io_in_from_accumu_mat_16(Quant_io_in_from_accumu_mat_16),
    .io_in_from_accumu_mat_17(Quant_io_in_from_accumu_mat_17),
    .io_in_from_accumu_mat_18(Quant_io_in_from_accumu_mat_18),
    .io_in_from_accumu_mat_19(Quant_io_in_from_accumu_mat_19),
    .io_in_from_accumu_mat_20(Quant_io_in_from_accumu_mat_20),
    .io_in_from_accumu_mat_21(Quant_io_in_from_accumu_mat_21),
    .io_in_from_accumu_mat_22(Quant_io_in_from_accumu_mat_22),
    .io_in_from_accumu_mat_23(Quant_io_in_from_accumu_mat_23),
    .io_in_from_accumu_mat_24(Quant_io_in_from_accumu_mat_24),
    .io_in_from_accumu_mat_25(Quant_io_in_from_accumu_mat_25),
    .io_in_from_accumu_mat_26(Quant_io_in_from_accumu_mat_26),
    .io_in_from_accumu_mat_27(Quant_io_in_from_accumu_mat_27),
    .io_in_from_accumu_mat_28(Quant_io_in_from_accumu_mat_28),
    .io_in_from_accumu_mat_29(Quant_io_in_from_accumu_mat_29),
    .io_in_from_accumu_mat_30(Quant_io_in_from_accumu_mat_30),
    .io_in_from_accumu_mat_31(Quant_io_in_from_accumu_mat_31),
    .io_in_from_accumu_mat_32(Quant_io_in_from_accumu_mat_32),
    .io_in_from_accumu_mat_33(Quant_io_in_from_accumu_mat_33),
    .io_in_from_accumu_mat_34(Quant_io_in_from_accumu_mat_34),
    .io_in_from_accumu_mat_35(Quant_io_in_from_accumu_mat_35),
    .io_in_from_accumu_mat_36(Quant_io_in_from_accumu_mat_36),
    .io_in_from_accumu_mat_37(Quant_io_in_from_accumu_mat_37),
    .io_in_from_accumu_mat_38(Quant_io_in_from_accumu_mat_38),
    .io_in_from_accumu_mat_39(Quant_io_in_from_accumu_mat_39),
    .io_in_from_accumu_mat_40(Quant_io_in_from_accumu_mat_40),
    .io_in_from_accumu_mat_41(Quant_io_in_from_accumu_mat_41),
    .io_in_from_accumu_mat_42(Quant_io_in_from_accumu_mat_42),
    .io_in_from_accumu_mat_43(Quant_io_in_from_accumu_mat_43),
    .io_in_from_accumu_mat_44(Quant_io_in_from_accumu_mat_44),
    .io_in_from_accumu_mat_45(Quant_io_in_from_accumu_mat_45),
    .io_in_from_accumu_mat_46(Quant_io_in_from_accumu_mat_46),
    .io_in_from_accumu_mat_47(Quant_io_in_from_accumu_mat_47),
    .io_in_from_accumu_mat_48(Quant_io_in_from_accumu_mat_48),
    .io_in_from_accumu_mat_49(Quant_io_in_from_accumu_mat_49),
    .io_in_from_accumu_mat_50(Quant_io_in_from_accumu_mat_50),
    .io_in_from_accumu_mat_51(Quant_io_in_from_accumu_mat_51),
    .io_in_from_accumu_mat_52(Quant_io_in_from_accumu_mat_52),
    .io_in_from_accumu_mat_53(Quant_io_in_from_accumu_mat_53),
    .io_in_from_accumu_mat_54(Quant_io_in_from_accumu_mat_54),
    .io_in_from_accumu_mat_55(Quant_io_in_from_accumu_mat_55),
    .io_in_from_accumu_mat_56(Quant_io_in_from_accumu_mat_56),
    .io_in_from_accumu_mat_57(Quant_io_in_from_accumu_mat_57),
    .io_in_from_accumu_mat_58(Quant_io_in_from_accumu_mat_58),
    .io_in_from_accumu_mat_59(Quant_io_in_from_accumu_mat_59),
    .io_in_from_accumu_mat_60(Quant_io_in_from_accumu_mat_60),
    .io_in_from_accumu_mat_61(Quant_io_in_from_accumu_mat_61),
    .io_in_from_accumu_mat_62(Quant_io_in_from_accumu_mat_62),
    .io_in_from_accumu_mat_63(Quant_io_in_from_accumu_mat_63),
    .io_result_mat_0(Quant_io_result_mat_0),
    .io_result_mat_1(Quant_io_result_mat_1),
    .io_result_mat_2(Quant_io_result_mat_2),
    .io_result_mat_3(Quant_io_result_mat_3),
    .io_result_mat_4(Quant_io_result_mat_4),
    .io_result_mat_5(Quant_io_result_mat_5),
    .io_result_mat_6(Quant_io_result_mat_6),
    .io_result_mat_7(Quant_io_result_mat_7),
    .io_result_mat_8(Quant_io_result_mat_8),
    .io_result_mat_9(Quant_io_result_mat_9),
    .io_result_mat_10(Quant_io_result_mat_10),
    .io_result_mat_11(Quant_io_result_mat_11),
    .io_result_mat_12(Quant_io_result_mat_12),
    .io_result_mat_13(Quant_io_result_mat_13),
    .io_result_mat_14(Quant_io_result_mat_14),
    .io_result_mat_15(Quant_io_result_mat_15),
    .io_result_mat_16(Quant_io_result_mat_16),
    .io_result_mat_17(Quant_io_result_mat_17),
    .io_result_mat_18(Quant_io_result_mat_18),
    .io_result_mat_19(Quant_io_result_mat_19),
    .io_result_mat_20(Quant_io_result_mat_20),
    .io_result_mat_21(Quant_io_result_mat_21),
    .io_result_mat_22(Quant_io_result_mat_22),
    .io_result_mat_23(Quant_io_result_mat_23),
    .io_result_mat_24(Quant_io_result_mat_24),
    .io_result_mat_25(Quant_io_result_mat_25),
    .io_result_mat_26(Quant_io_result_mat_26),
    .io_result_mat_27(Quant_io_result_mat_27),
    .io_result_mat_28(Quant_io_result_mat_28),
    .io_result_mat_29(Quant_io_result_mat_29),
    .io_result_mat_30(Quant_io_result_mat_30),
    .io_result_mat_31(Quant_io_result_mat_31),
    .io_result_mat_32(Quant_io_result_mat_32),
    .io_result_mat_33(Quant_io_result_mat_33),
    .io_result_mat_34(Quant_io_result_mat_34),
    .io_result_mat_35(Quant_io_result_mat_35),
    .io_result_mat_36(Quant_io_result_mat_36),
    .io_result_mat_37(Quant_io_result_mat_37),
    .io_result_mat_38(Quant_io_result_mat_38),
    .io_result_mat_39(Quant_io_result_mat_39),
    .io_result_mat_40(Quant_io_result_mat_40),
    .io_result_mat_41(Quant_io_result_mat_41),
    .io_result_mat_42(Quant_io_result_mat_42),
    .io_result_mat_43(Quant_io_result_mat_43),
    .io_result_mat_44(Quant_io_result_mat_44),
    .io_result_mat_45(Quant_io_result_mat_45),
    .io_result_mat_46(Quant_io_result_mat_46),
    .io_result_mat_47(Quant_io_result_mat_47),
    .io_result_mat_48(Quant_io_result_mat_48),
    .io_result_mat_49(Quant_io_result_mat_49),
    .io_result_mat_50(Quant_io_result_mat_50),
    .io_result_mat_51(Quant_io_result_mat_51),
    .io_result_mat_52(Quant_io_result_mat_52),
    .io_result_mat_53(Quant_io_result_mat_53),
    .io_result_mat_54(Quant_io_result_mat_54),
    .io_result_mat_55(Quant_io_result_mat_55),
    .io_result_mat_56(Quant_io_result_mat_56),
    .io_result_mat_57(Quant_io_result_mat_57),
    .io_result_mat_58(Quant_io_result_mat_58),
    .io_result_mat_59(Quant_io_result_mat_59),
    .io_result_mat_60(Quant_io_result_mat_60),
    .io_result_mat_61(Quant_io_result_mat_61),
    .io_result_mat_62(Quant_io_result_mat_62),
    .io_result_mat_63(Quant_io_result_mat_63),
    .io_quant_in_in_q(Quant_io_quant_in_in_q),
    .io_quant_in_out_q(Quant_io_quant_in_out_q)
  );
  WriteSwitch WriteSwitch ( // @[top.scala 22:30]
    .io_valid_in_0(WriteSwitch_io_valid_in_0),
    .io_valid_out(WriteSwitch_io_valid_out),
    .io_input_0_mat_0(WriteSwitch_io_input_0_mat_0),
    .io_input_0_mat_1(WriteSwitch_io_input_0_mat_1),
    .io_input_0_mat_2(WriteSwitch_io_input_0_mat_2),
    .io_input_0_mat_3(WriteSwitch_io_input_0_mat_3),
    .io_input_0_mat_4(WriteSwitch_io_input_0_mat_4),
    .io_input_0_mat_5(WriteSwitch_io_input_0_mat_5),
    .io_input_0_mat_6(WriteSwitch_io_input_0_mat_6),
    .io_input_0_mat_7(WriteSwitch_io_input_0_mat_7),
    .io_input_0_mat_8(WriteSwitch_io_input_0_mat_8),
    .io_input_0_mat_9(WriteSwitch_io_input_0_mat_9),
    .io_input_0_mat_10(WriteSwitch_io_input_0_mat_10),
    .io_input_0_mat_11(WriteSwitch_io_input_0_mat_11),
    .io_input_0_mat_12(WriteSwitch_io_input_0_mat_12),
    .io_input_0_mat_13(WriteSwitch_io_input_0_mat_13),
    .io_input_0_mat_14(WriteSwitch_io_input_0_mat_14),
    .io_input_0_mat_15(WriteSwitch_io_input_0_mat_15),
    .io_input_0_mat_16(WriteSwitch_io_input_0_mat_16),
    .io_input_0_mat_17(WriteSwitch_io_input_0_mat_17),
    .io_input_0_mat_18(WriteSwitch_io_input_0_mat_18),
    .io_input_0_mat_19(WriteSwitch_io_input_0_mat_19),
    .io_input_0_mat_20(WriteSwitch_io_input_0_mat_20),
    .io_input_0_mat_21(WriteSwitch_io_input_0_mat_21),
    .io_input_0_mat_22(WriteSwitch_io_input_0_mat_22),
    .io_input_0_mat_23(WriteSwitch_io_input_0_mat_23),
    .io_input_0_mat_24(WriteSwitch_io_input_0_mat_24),
    .io_input_0_mat_25(WriteSwitch_io_input_0_mat_25),
    .io_input_0_mat_26(WriteSwitch_io_input_0_mat_26),
    .io_input_0_mat_27(WriteSwitch_io_input_0_mat_27),
    .io_input_0_mat_28(WriteSwitch_io_input_0_mat_28),
    .io_input_0_mat_29(WriteSwitch_io_input_0_mat_29),
    .io_input_0_mat_30(WriteSwitch_io_input_0_mat_30),
    .io_input_0_mat_31(WriteSwitch_io_input_0_mat_31),
    .io_input_0_mat_32(WriteSwitch_io_input_0_mat_32),
    .io_input_0_mat_33(WriteSwitch_io_input_0_mat_33),
    .io_input_0_mat_34(WriteSwitch_io_input_0_mat_34),
    .io_input_0_mat_35(WriteSwitch_io_input_0_mat_35),
    .io_input_0_mat_36(WriteSwitch_io_input_0_mat_36),
    .io_input_0_mat_37(WriteSwitch_io_input_0_mat_37),
    .io_input_0_mat_38(WriteSwitch_io_input_0_mat_38),
    .io_input_0_mat_39(WriteSwitch_io_input_0_mat_39),
    .io_input_0_mat_40(WriteSwitch_io_input_0_mat_40),
    .io_input_0_mat_41(WriteSwitch_io_input_0_mat_41),
    .io_input_0_mat_42(WriteSwitch_io_input_0_mat_42),
    .io_input_0_mat_43(WriteSwitch_io_input_0_mat_43),
    .io_input_0_mat_44(WriteSwitch_io_input_0_mat_44),
    .io_input_0_mat_45(WriteSwitch_io_input_0_mat_45),
    .io_input_0_mat_46(WriteSwitch_io_input_0_mat_46),
    .io_input_0_mat_47(WriteSwitch_io_input_0_mat_47),
    .io_input_0_mat_48(WriteSwitch_io_input_0_mat_48),
    .io_input_0_mat_49(WriteSwitch_io_input_0_mat_49),
    .io_input_0_mat_50(WriteSwitch_io_input_0_mat_50),
    .io_input_0_mat_51(WriteSwitch_io_input_0_mat_51),
    .io_input_0_mat_52(WriteSwitch_io_input_0_mat_52),
    .io_input_0_mat_53(WriteSwitch_io_input_0_mat_53),
    .io_input_0_mat_54(WriteSwitch_io_input_0_mat_54),
    .io_input_0_mat_55(WriteSwitch_io_input_0_mat_55),
    .io_input_0_mat_56(WriteSwitch_io_input_0_mat_56),
    .io_input_0_mat_57(WriteSwitch_io_input_0_mat_57),
    .io_input_0_mat_58(WriteSwitch_io_input_0_mat_58),
    .io_input_0_mat_59(WriteSwitch_io_input_0_mat_59),
    .io_input_0_mat_60(WriteSwitch_io_input_0_mat_60),
    .io_input_0_mat_61(WriteSwitch_io_input_0_mat_61),
    .io_input_0_mat_62(WriteSwitch_io_input_0_mat_62),
    .io_input_0_mat_63(WriteSwitch_io_input_0_mat_63),
    .io_output_mat_0(WriteSwitch_io_output_mat_0),
    .io_output_mat_1(WriteSwitch_io_output_mat_1),
    .io_output_mat_2(WriteSwitch_io_output_mat_2),
    .io_output_mat_3(WriteSwitch_io_output_mat_3),
    .io_output_mat_4(WriteSwitch_io_output_mat_4),
    .io_output_mat_5(WriteSwitch_io_output_mat_5),
    .io_output_mat_6(WriteSwitch_io_output_mat_6),
    .io_output_mat_7(WriteSwitch_io_output_mat_7),
    .io_output_mat_8(WriteSwitch_io_output_mat_8),
    .io_output_mat_9(WriteSwitch_io_output_mat_9),
    .io_output_mat_10(WriteSwitch_io_output_mat_10),
    .io_output_mat_11(WriteSwitch_io_output_mat_11),
    .io_output_mat_12(WriteSwitch_io_output_mat_12),
    .io_output_mat_13(WriteSwitch_io_output_mat_13),
    .io_output_mat_14(WriteSwitch_io_output_mat_14),
    .io_output_mat_15(WriteSwitch_io_output_mat_15),
    .io_output_mat_16(WriteSwitch_io_output_mat_16),
    .io_output_mat_17(WriteSwitch_io_output_mat_17),
    .io_output_mat_18(WriteSwitch_io_output_mat_18),
    .io_output_mat_19(WriteSwitch_io_output_mat_19),
    .io_output_mat_20(WriteSwitch_io_output_mat_20),
    .io_output_mat_21(WriteSwitch_io_output_mat_21),
    .io_output_mat_22(WriteSwitch_io_output_mat_22),
    .io_output_mat_23(WriteSwitch_io_output_mat_23),
    .io_output_mat_24(WriteSwitch_io_output_mat_24),
    .io_output_mat_25(WriteSwitch_io_output_mat_25),
    .io_output_mat_26(WriteSwitch_io_output_mat_26),
    .io_output_mat_27(WriteSwitch_io_output_mat_27),
    .io_output_mat_28(WriteSwitch_io_output_mat_28),
    .io_output_mat_29(WriteSwitch_io_output_mat_29),
    .io_output_mat_30(WriteSwitch_io_output_mat_30),
    .io_output_mat_31(WriteSwitch_io_output_mat_31),
    .io_output_mat_32(WriteSwitch_io_output_mat_32),
    .io_output_mat_33(WriteSwitch_io_output_mat_33),
    .io_output_mat_34(WriteSwitch_io_output_mat_34),
    .io_output_mat_35(WriteSwitch_io_output_mat_35),
    .io_output_mat_36(WriteSwitch_io_output_mat_36),
    .io_output_mat_37(WriteSwitch_io_output_mat_37),
    .io_output_mat_38(WriteSwitch_io_output_mat_38),
    .io_output_mat_39(WriteSwitch_io_output_mat_39),
    .io_output_mat_40(WriteSwitch_io_output_mat_40),
    .io_output_mat_41(WriteSwitch_io_output_mat_41),
    .io_output_mat_42(WriteSwitch_io_output_mat_42),
    .io_output_mat_43(WriteSwitch_io_output_mat_43),
    .io_output_mat_44(WriteSwitch_io_output_mat_44),
    .io_output_mat_45(WriteSwitch_io_output_mat_45),
    .io_output_mat_46(WriteSwitch_io_output_mat_46),
    .io_output_mat_47(WriteSwitch_io_output_mat_47),
    .io_output_mat_48(WriteSwitch_io_output_mat_48),
    .io_output_mat_49(WriteSwitch_io_output_mat_49),
    .io_output_mat_50(WriteSwitch_io_output_mat_50),
    .io_output_mat_51(WriteSwitch_io_output_mat_51),
    .io_output_mat_52(WriteSwitch_io_output_mat_52),
    .io_output_mat_53(WriteSwitch_io_output_mat_53),
    .io_output_mat_54(WriteSwitch_io_output_mat_54),
    .io_output_mat_55(WriteSwitch_io_output_mat_55),
    .io_output_mat_56(WriteSwitch_io_output_mat_56),
    .io_output_mat_57(WriteSwitch_io_output_mat_57),
    .io_output_mat_58(WriteSwitch_io_output_mat_58),
    .io_output_mat_59(WriteSwitch_io_output_mat_59),
    .io_output_mat_60(WriteSwitch_io_output_mat_60),
    .io_output_mat_61(WriteSwitch_io_output_mat_61),
    .io_output_mat_62(WriteSwitch_io_output_mat_62),
    .io_output_mat_63(WriteSwitch_io_output_mat_63)
  );
  RealWriter RealWriter ( // @[top.scala 23:24]
    .clock(RealWriter_clock),
    .reset(RealWriter_reset),
    .io_valid_in(RealWriter_io_valid_in),
    .io_valid_out(RealWriter_io_valid_out),
    .io_flag_job(RealWriter_io_flag_job),
    .io_in_from_quant_mat_0(RealWriter_io_in_from_quant_mat_0),
    .io_in_from_quant_mat_1(RealWriter_io_in_from_quant_mat_1),
    .io_in_from_quant_mat_2(RealWriter_io_in_from_quant_mat_2),
    .io_in_from_quant_mat_3(RealWriter_io_in_from_quant_mat_3),
    .io_in_from_quant_mat_4(RealWriter_io_in_from_quant_mat_4),
    .io_in_from_quant_mat_5(RealWriter_io_in_from_quant_mat_5),
    .io_in_from_quant_mat_6(RealWriter_io_in_from_quant_mat_6),
    .io_in_from_quant_mat_7(RealWriter_io_in_from_quant_mat_7),
    .io_in_from_quant_mat_8(RealWriter_io_in_from_quant_mat_8),
    .io_in_from_quant_mat_9(RealWriter_io_in_from_quant_mat_9),
    .io_in_from_quant_mat_10(RealWriter_io_in_from_quant_mat_10),
    .io_in_from_quant_mat_11(RealWriter_io_in_from_quant_mat_11),
    .io_in_from_quant_mat_12(RealWriter_io_in_from_quant_mat_12),
    .io_in_from_quant_mat_13(RealWriter_io_in_from_quant_mat_13),
    .io_in_from_quant_mat_14(RealWriter_io_in_from_quant_mat_14),
    .io_in_from_quant_mat_15(RealWriter_io_in_from_quant_mat_15),
    .io_in_from_quant_mat_16(RealWriter_io_in_from_quant_mat_16),
    .io_in_from_quant_mat_17(RealWriter_io_in_from_quant_mat_17),
    .io_in_from_quant_mat_18(RealWriter_io_in_from_quant_mat_18),
    .io_in_from_quant_mat_19(RealWriter_io_in_from_quant_mat_19),
    .io_in_from_quant_mat_20(RealWriter_io_in_from_quant_mat_20),
    .io_in_from_quant_mat_21(RealWriter_io_in_from_quant_mat_21),
    .io_in_from_quant_mat_22(RealWriter_io_in_from_quant_mat_22),
    .io_in_from_quant_mat_23(RealWriter_io_in_from_quant_mat_23),
    .io_in_from_quant_mat_24(RealWriter_io_in_from_quant_mat_24),
    .io_in_from_quant_mat_25(RealWriter_io_in_from_quant_mat_25),
    .io_in_from_quant_mat_26(RealWriter_io_in_from_quant_mat_26),
    .io_in_from_quant_mat_27(RealWriter_io_in_from_quant_mat_27),
    .io_in_from_quant_mat_28(RealWriter_io_in_from_quant_mat_28),
    .io_in_from_quant_mat_29(RealWriter_io_in_from_quant_mat_29),
    .io_in_from_quant_mat_30(RealWriter_io_in_from_quant_mat_30),
    .io_in_from_quant_mat_31(RealWriter_io_in_from_quant_mat_31),
    .io_in_from_quant_mat_32(RealWriter_io_in_from_quant_mat_32),
    .io_in_from_quant_mat_33(RealWriter_io_in_from_quant_mat_33),
    .io_in_from_quant_mat_34(RealWriter_io_in_from_quant_mat_34),
    .io_in_from_quant_mat_35(RealWriter_io_in_from_quant_mat_35),
    .io_in_from_quant_mat_36(RealWriter_io_in_from_quant_mat_36),
    .io_in_from_quant_mat_37(RealWriter_io_in_from_quant_mat_37),
    .io_in_from_quant_mat_38(RealWriter_io_in_from_quant_mat_38),
    .io_in_from_quant_mat_39(RealWriter_io_in_from_quant_mat_39),
    .io_in_from_quant_mat_40(RealWriter_io_in_from_quant_mat_40),
    .io_in_from_quant_mat_41(RealWriter_io_in_from_quant_mat_41),
    .io_in_from_quant_mat_42(RealWriter_io_in_from_quant_mat_42),
    .io_in_from_quant_mat_43(RealWriter_io_in_from_quant_mat_43),
    .io_in_from_quant_mat_44(RealWriter_io_in_from_quant_mat_44),
    .io_in_from_quant_mat_45(RealWriter_io_in_from_quant_mat_45),
    .io_in_from_quant_mat_46(RealWriter_io_in_from_quant_mat_46),
    .io_in_from_quant_mat_47(RealWriter_io_in_from_quant_mat_47),
    .io_in_from_quant_mat_48(RealWriter_io_in_from_quant_mat_48),
    .io_in_from_quant_mat_49(RealWriter_io_in_from_quant_mat_49),
    .io_in_from_quant_mat_50(RealWriter_io_in_from_quant_mat_50),
    .io_in_from_quant_mat_51(RealWriter_io_in_from_quant_mat_51),
    .io_in_from_quant_mat_52(RealWriter_io_in_from_quant_mat_52),
    .io_in_from_quant_mat_53(RealWriter_io_in_from_quant_mat_53),
    .io_in_from_quant_mat_54(RealWriter_io_in_from_quant_mat_54),
    .io_in_from_quant_mat_55(RealWriter_io_in_from_quant_mat_55),
    .io_in_from_quant_mat_56(RealWriter_io_in_from_quant_mat_56),
    .io_in_from_quant_mat_57(RealWriter_io_in_from_quant_mat_57),
    .io_in_from_quant_mat_58(RealWriter_io_in_from_quant_mat_58),
    .io_in_from_quant_mat_59(RealWriter_io_in_from_quant_mat_59),
    .io_in_from_quant_mat_60(RealWriter_io_in_from_quant_mat_60),
    .io_in_from_quant_mat_61(RealWriter_io_in_from_quant_mat_61),
    .io_in_from_quant_mat_62(RealWriter_io_in_from_quant_mat_62),
    .io_in_from_quant_mat_63(RealWriter_io_in_from_quant_mat_63),
    .io_job_job_0_big_begin_addr(RealWriter_io_job_job_0_big_begin_addr),
    .io_job_job_0_big_max_addr(RealWriter_io_job_job_0_big_max_addr),
    .io_job_job_0_big_cnt_ic_end(RealWriter_io_job_job_0_big_cnt_ic_end),
    .io_job_job_0_big_a(RealWriter_io_job_job_0_big_a),
    .io_job_job_0_small_0_begin_addr(RealWriter_io_job_job_0_small_0_begin_addr),
    .io_job_job_0_small_0_max_addr(RealWriter_io_job_job_0_small_0_max_addr),
    .io_job_job_0_small_0_cnt_y_end(RealWriter_io_job_job_0_small_0_cnt_y_end),
    .io_job_job_0_small_0_cnt_ic_end(RealWriter_io_job_job_0_small_0_cnt_ic_end),
    .io_job_job_0_small_0_a(RealWriter_io_job_job_0_small_0_a),
    .io_job_job_0_small_0_ano_bank_id(RealWriter_io_job_job_0_small_0_ano_bank_id),
    .io_job_job_0_small_1_begin_addr(RealWriter_io_job_job_0_small_1_begin_addr),
    .io_job_job_0_small_1_max_addr(RealWriter_io_job_job_0_small_1_max_addr),
    .io_job_job_0_small_1_bank_id(RealWriter_io_job_job_0_small_1_bank_id),
    .io_job_job_0_small_1_cnt_y_end(RealWriter_io_job_job_0_small_1_cnt_y_end),
    .io_job_job_0_small_1_cnt_ic_end(RealWriter_io_job_job_0_small_1_cnt_ic_end),
    .io_job_job_0_small_1_a(RealWriter_io_job_job_0_small_1_a),
    .io_job_job_0_small_1_ano_bank_id(RealWriter_io_job_job_0_small_1_ano_bank_id),
    .io_job_job_1_big_begin_addr(RealWriter_io_job_job_1_big_begin_addr),
    .io_job_job_1_big_max_addr(RealWriter_io_job_job_1_big_max_addr),
    .io_job_job_1_big_bank_id(RealWriter_io_job_job_1_big_bank_id),
    .io_job_job_1_big_cnt_ic_end(RealWriter_io_job_job_1_big_cnt_ic_end),
    .io_job_job_1_big_a(RealWriter_io_job_job_1_big_a),
    .io_job_job_1_small_0_begin_addr(RealWriter_io_job_job_1_small_0_begin_addr),
    .io_job_job_1_small_0_max_addr(RealWriter_io_job_job_1_small_0_max_addr),
    .io_job_job_1_small_0_bank_id(RealWriter_io_job_job_1_small_0_bank_id),
    .io_job_job_1_small_0_cnt_y_end(RealWriter_io_job_job_1_small_0_cnt_y_end),
    .io_job_job_1_small_0_cnt_ic_end(RealWriter_io_job_job_1_small_0_cnt_ic_end),
    .io_job_job_1_small_0_a(RealWriter_io_job_job_1_small_0_a),
    .io_job_job_1_small_0_ano_bank_id(RealWriter_io_job_job_1_small_0_ano_bank_id),
    .io_job_job_1_small_1_begin_addr(RealWriter_io_job_job_1_small_1_begin_addr),
    .io_job_job_1_small_1_max_addr(RealWriter_io_job_job_1_small_1_max_addr),
    .io_job_job_1_small_1_bank_id(RealWriter_io_job_job_1_small_1_bank_id),
    .io_job_job_1_small_1_cnt_y_end(RealWriter_io_job_job_1_small_1_cnt_y_end),
    .io_job_job_1_small_1_cnt_ic_end(RealWriter_io_job_job_1_small_1_cnt_ic_end),
    .io_job_job_1_small_1_a(RealWriter_io_job_job_1_small_1_a),
    .io_job_job_1_small_1_ano_bank_id(RealWriter_io_job_job_1_small_1_ano_bank_id),
    .io_job_out_chan(RealWriter_io_job_out_chan),
    .io_to_bigbank_data_0(RealWriter_io_to_bigbank_data_0),
    .io_to_bigbank_data_1(RealWriter_io_to_bigbank_data_1),
    .io_to_bigbank_data_2(RealWriter_io_to_bigbank_data_2),
    .io_to_bigbank_data_3(RealWriter_io_to_bigbank_data_3),
    .io_to_bigbank_data_4(RealWriter_io_to_bigbank_data_4),
    .io_to_bigbank_data_5(RealWriter_io_to_bigbank_data_5),
    .io_to_bigbank_data_6(RealWriter_io_to_bigbank_data_6),
    .io_to_bigbank_data_7(RealWriter_io_to_bigbank_data_7),
    .io_to_bigbank_data_8(RealWriter_io_to_bigbank_data_8),
    .io_to_bigbank_data_9(RealWriter_io_to_bigbank_data_9),
    .io_to_bigbank_data_10(RealWriter_io_to_bigbank_data_10),
    .io_to_bigbank_data_11(RealWriter_io_to_bigbank_data_11),
    .io_to_bigbank_data_12(RealWriter_io_to_bigbank_data_12),
    .io_to_bigbank_data_13(RealWriter_io_to_bigbank_data_13),
    .io_to_bigbank_data_14(RealWriter_io_to_bigbank_data_14),
    .io_to_bigbank_data_15(RealWriter_io_to_bigbank_data_15),
    .io_to_bigbank_data_16(RealWriter_io_to_bigbank_data_16),
    .io_to_bigbank_data_17(RealWriter_io_to_bigbank_data_17),
    .io_to_bigbank_data_18(RealWriter_io_to_bigbank_data_18),
    .io_to_bigbank_data_19(RealWriter_io_to_bigbank_data_19),
    .io_to_bigbank_data_20(RealWriter_io_to_bigbank_data_20),
    .io_to_bigbank_data_21(RealWriter_io_to_bigbank_data_21),
    .io_to_bigbank_data_22(RealWriter_io_to_bigbank_data_22),
    .io_to_bigbank_data_23(RealWriter_io_to_bigbank_data_23),
    .io_to_bigbank_data_24(RealWriter_io_to_bigbank_data_24),
    .io_to_bigbank_data_25(RealWriter_io_to_bigbank_data_25),
    .io_to_bigbank_data_26(RealWriter_io_to_bigbank_data_26),
    .io_to_bigbank_data_27(RealWriter_io_to_bigbank_data_27),
    .io_to_bigbank_data_28(RealWriter_io_to_bigbank_data_28),
    .io_to_bigbank_data_29(RealWriter_io_to_bigbank_data_29),
    .io_to_bigbank_data_30(RealWriter_io_to_bigbank_data_30),
    .io_to_bigbank_data_31(RealWriter_io_to_bigbank_data_31),
    .io_to_bigbank_data_32(RealWriter_io_to_bigbank_data_32),
    .io_to_bigbank_data_33(RealWriter_io_to_bigbank_data_33),
    .io_to_bigbank_data_34(RealWriter_io_to_bigbank_data_34),
    .io_to_bigbank_data_35(RealWriter_io_to_bigbank_data_35),
    .io_to_bigbank_data_36(RealWriter_io_to_bigbank_data_36),
    .io_to_bigbank_data_37(RealWriter_io_to_bigbank_data_37),
    .io_to_bigbank_data_38(RealWriter_io_to_bigbank_data_38),
    .io_to_bigbank_data_39(RealWriter_io_to_bigbank_data_39),
    .io_to_bigbank_data_40(RealWriter_io_to_bigbank_data_40),
    .io_to_bigbank_data_41(RealWriter_io_to_bigbank_data_41),
    .io_to_bigbank_data_42(RealWriter_io_to_bigbank_data_42),
    .io_to_bigbank_data_43(RealWriter_io_to_bigbank_data_43),
    .io_to_bigbank_data_44(RealWriter_io_to_bigbank_data_44),
    .io_to_bigbank_data_45(RealWriter_io_to_bigbank_data_45),
    .io_to_bigbank_data_46(RealWriter_io_to_bigbank_data_46),
    .io_to_bigbank_data_47(RealWriter_io_to_bigbank_data_47),
    .io_to_smallbank_0_data_0(RealWriter_io_to_smallbank_0_data_0),
    .io_to_smallbank_0_data_1(RealWriter_io_to_smallbank_0_data_1),
    .io_to_smallbank_0_data_2(RealWriter_io_to_smallbank_0_data_2),
    .io_to_smallbank_0_data_3(RealWriter_io_to_smallbank_0_data_3),
    .io_to_smallbank_0_data_4(RealWriter_io_to_smallbank_0_data_4),
    .io_to_smallbank_0_data_5(RealWriter_io_to_smallbank_0_data_5),
    .io_to_smallbank_0_data_6(RealWriter_io_to_smallbank_0_data_6),
    .io_to_smallbank_0_data_7(RealWriter_io_to_smallbank_0_data_7),
    .io_to_smallbank_1_data_0(RealWriter_io_to_smallbank_1_data_0),
    .io_to_smallbank_1_data_1(RealWriter_io_to_smallbank_1_data_1),
    .io_to_smallbank_1_data_2(RealWriter_io_to_smallbank_1_data_2),
    .io_to_smallbank_1_data_3(RealWriter_io_to_smallbank_1_data_3),
    .io_to_smallbank_1_data_4(RealWriter_io_to_smallbank_1_data_4),
    .io_to_smallbank_1_data_5(RealWriter_io_to_smallbank_1_data_5),
    .io_to_smallbank_1_data_6(RealWriter_io_to_smallbank_1_data_6),
    .io_to_smallbank_1_data_7(RealWriter_io_to_smallbank_1_data_7),
    .io_to_banks_addrs_0_addr(RealWriter_io_to_banks_addrs_0_addr),
    .io_to_banks_addrs_0_bank_id(RealWriter_io_to_banks_addrs_0_bank_id),
    .io_to_banks_addrs_1_addr(RealWriter_io_to_banks_addrs_1_addr),
    .io_to_banks_addrs_1_bank_id(RealWriter_io_to_banks_addrs_1_bank_id),
    .io_to_banks_addrs_2_addr(RealWriter_io_to_banks_addrs_2_addr),
    .io_to_banks_addrs_2_bank_id(RealWriter_io_to_banks_addrs_2_bank_id)
  );
  ROMWeight ROMWeight ( // @[top.scala 26:28]
    .clock(ROMWeight_clock),
    .io_addr(ROMWeight_io_addr),
    .io_out_0(ROMWeight_io_out_0),
    .io_out_1(ROMWeight_io_out_1),
    .io_out_2(ROMWeight_io_out_2),
    .io_out_3(ROMWeight_io_out_3),
    .io_out_4(ROMWeight_io_out_4),
    .io_out_5(ROMWeight_io_out_5),
    .io_out_6(ROMWeight_io_out_6),
    .io_out_7(ROMWeight_io_out_7),
    .io_out_8(ROMWeight_io_out_8)
  );
  ROMBias ROMBias ( // @[top.scala 27:26]
    .clock(ROMBias_clock),
    .io_addr(ROMBias_io_addr),
    .io_out(ROMBias_io_out)
  );
  RAMGroup RAMGroup ( // @[top.scala 28:22]
    .clock(RAMGroup_clock),
    .reset(RAMGroup_reset),
    .io_rd_valid_in(RAMGroup_io_rd_valid_in),
    .io_rd_valid_out(RAMGroup_io_rd_valid_out),
    .io_rd_addr1_addrs_0_bank_id(RAMGroup_io_rd_addr1_addrs_0_bank_id),
    .io_rd_addr1_addrs_1_addr(RAMGroup_io_rd_addr1_addrs_1_addr),
    .io_rd_addr2_addrs_1_addr(RAMGroup_io_rd_addr2_addrs_1_addr),
    .io_rd_big_0_data_0(RAMGroup_io_rd_big_0_data_0),
    .io_rd_big_0_data_1(RAMGroup_io_rd_big_0_data_1),
    .io_rd_big_0_data_2(RAMGroup_io_rd_big_0_data_2),
    .io_rd_big_0_data_3(RAMGroup_io_rd_big_0_data_3),
    .io_rd_big_0_data_4(RAMGroup_io_rd_big_0_data_4),
    .io_rd_big_0_data_5(RAMGroup_io_rd_big_0_data_5),
    .io_rd_big_0_data_6(RAMGroup_io_rd_big_0_data_6),
    .io_rd_big_0_data_7(RAMGroup_io_rd_big_0_data_7),
    .io_rd_big_0_data_8(RAMGroup_io_rd_big_0_data_8),
    .io_rd_big_0_data_9(RAMGroup_io_rd_big_0_data_9),
    .io_rd_big_0_data_10(RAMGroup_io_rd_big_0_data_10),
    .io_rd_big_0_data_11(RAMGroup_io_rd_big_0_data_11),
    .io_rd_big_0_data_12(RAMGroup_io_rd_big_0_data_12),
    .io_rd_big_0_data_13(RAMGroup_io_rd_big_0_data_13),
    .io_rd_big_0_data_14(RAMGroup_io_rd_big_0_data_14),
    .io_rd_big_0_data_15(RAMGroup_io_rd_big_0_data_15),
    .io_rd_big_0_data_16(RAMGroup_io_rd_big_0_data_16),
    .io_rd_big_0_data_17(RAMGroup_io_rd_big_0_data_17),
    .io_rd_big_0_data_18(RAMGroup_io_rd_big_0_data_18),
    .io_rd_big_0_data_19(RAMGroup_io_rd_big_0_data_19),
    .io_rd_big_0_data_20(RAMGroup_io_rd_big_0_data_20),
    .io_rd_big_0_data_21(RAMGroup_io_rd_big_0_data_21),
    .io_rd_big_0_data_22(RAMGroup_io_rd_big_0_data_22),
    .io_rd_big_0_data_23(RAMGroup_io_rd_big_0_data_23),
    .io_rd_big_0_data_24(RAMGroup_io_rd_big_0_data_24),
    .io_rd_big_0_data_25(RAMGroup_io_rd_big_0_data_25),
    .io_rd_big_0_data_26(RAMGroup_io_rd_big_0_data_26),
    .io_rd_big_0_data_27(RAMGroup_io_rd_big_0_data_27),
    .io_rd_big_0_data_28(RAMGroup_io_rd_big_0_data_28),
    .io_rd_big_0_data_29(RAMGroup_io_rd_big_0_data_29),
    .io_rd_big_0_data_30(RAMGroup_io_rd_big_0_data_30),
    .io_rd_big_0_data_31(RAMGroup_io_rd_big_0_data_31),
    .io_rd_big_0_data_32(RAMGroup_io_rd_big_0_data_32),
    .io_rd_big_0_data_33(RAMGroup_io_rd_big_0_data_33),
    .io_rd_big_0_data_34(RAMGroup_io_rd_big_0_data_34),
    .io_rd_big_0_data_35(RAMGroup_io_rd_big_0_data_35),
    .io_rd_big_0_data_36(RAMGroup_io_rd_big_0_data_36),
    .io_rd_big_0_data_37(RAMGroup_io_rd_big_0_data_37),
    .io_rd_big_0_data_38(RAMGroup_io_rd_big_0_data_38),
    .io_rd_big_0_data_39(RAMGroup_io_rd_big_0_data_39),
    .io_rd_big_0_data_40(RAMGroup_io_rd_big_0_data_40),
    .io_rd_big_0_data_41(RAMGroup_io_rd_big_0_data_41),
    .io_rd_big_0_data_42(RAMGroup_io_rd_big_0_data_42),
    .io_rd_big_0_data_43(RAMGroup_io_rd_big_0_data_43),
    .io_rd_big_0_data_44(RAMGroup_io_rd_big_0_data_44),
    .io_rd_big_0_data_45(RAMGroup_io_rd_big_0_data_45),
    .io_rd_big_0_data_46(RAMGroup_io_rd_big_0_data_46),
    .io_rd_big_0_data_47(RAMGroup_io_rd_big_0_data_47),
    .io_rd_big_1_data_0(RAMGroup_io_rd_big_1_data_0),
    .io_rd_big_1_data_1(RAMGroup_io_rd_big_1_data_1),
    .io_rd_big_1_data_2(RAMGroup_io_rd_big_1_data_2),
    .io_rd_big_1_data_3(RAMGroup_io_rd_big_1_data_3),
    .io_rd_big_1_data_4(RAMGroup_io_rd_big_1_data_4),
    .io_rd_big_1_data_5(RAMGroup_io_rd_big_1_data_5),
    .io_rd_big_1_data_6(RAMGroup_io_rd_big_1_data_6),
    .io_rd_big_1_data_7(RAMGroup_io_rd_big_1_data_7),
    .io_rd_big_1_data_8(RAMGroup_io_rd_big_1_data_8),
    .io_rd_big_1_data_9(RAMGroup_io_rd_big_1_data_9),
    .io_rd_big_1_data_10(RAMGroup_io_rd_big_1_data_10),
    .io_rd_big_1_data_11(RAMGroup_io_rd_big_1_data_11),
    .io_rd_big_1_data_12(RAMGroup_io_rd_big_1_data_12),
    .io_rd_big_1_data_13(RAMGroup_io_rd_big_1_data_13),
    .io_rd_big_1_data_14(RAMGroup_io_rd_big_1_data_14),
    .io_rd_big_1_data_15(RAMGroup_io_rd_big_1_data_15),
    .io_rd_big_1_data_16(RAMGroup_io_rd_big_1_data_16),
    .io_rd_big_1_data_17(RAMGroup_io_rd_big_1_data_17),
    .io_rd_big_1_data_18(RAMGroup_io_rd_big_1_data_18),
    .io_rd_big_1_data_19(RAMGroup_io_rd_big_1_data_19),
    .io_rd_big_1_data_20(RAMGroup_io_rd_big_1_data_20),
    .io_rd_big_1_data_21(RAMGroup_io_rd_big_1_data_21),
    .io_rd_big_1_data_22(RAMGroup_io_rd_big_1_data_22),
    .io_rd_big_1_data_23(RAMGroup_io_rd_big_1_data_23),
    .io_rd_big_1_data_24(RAMGroup_io_rd_big_1_data_24),
    .io_rd_big_1_data_25(RAMGroup_io_rd_big_1_data_25),
    .io_rd_big_1_data_26(RAMGroup_io_rd_big_1_data_26),
    .io_rd_big_1_data_27(RAMGroup_io_rd_big_1_data_27),
    .io_rd_big_1_data_28(RAMGroup_io_rd_big_1_data_28),
    .io_rd_big_1_data_29(RAMGroup_io_rd_big_1_data_29),
    .io_rd_big_1_data_30(RAMGroup_io_rd_big_1_data_30),
    .io_rd_big_1_data_31(RAMGroup_io_rd_big_1_data_31),
    .io_rd_big_1_data_32(RAMGroup_io_rd_big_1_data_32),
    .io_rd_big_1_data_33(RAMGroup_io_rd_big_1_data_33),
    .io_rd_big_1_data_34(RAMGroup_io_rd_big_1_data_34),
    .io_rd_big_1_data_35(RAMGroup_io_rd_big_1_data_35),
    .io_rd_big_1_data_36(RAMGroup_io_rd_big_1_data_36),
    .io_rd_big_1_data_37(RAMGroup_io_rd_big_1_data_37),
    .io_rd_big_1_data_38(RAMGroup_io_rd_big_1_data_38),
    .io_rd_big_1_data_39(RAMGroup_io_rd_big_1_data_39),
    .io_rd_big_1_data_40(RAMGroup_io_rd_big_1_data_40),
    .io_rd_big_1_data_41(RAMGroup_io_rd_big_1_data_41),
    .io_rd_big_1_data_42(RAMGroup_io_rd_big_1_data_42),
    .io_rd_big_1_data_43(RAMGroup_io_rd_big_1_data_43),
    .io_rd_big_1_data_44(RAMGroup_io_rd_big_1_data_44),
    .io_rd_big_1_data_45(RAMGroup_io_rd_big_1_data_45),
    .io_rd_big_1_data_46(RAMGroup_io_rd_big_1_data_46),
    .io_rd_big_1_data_47(RAMGroup_io_rd_big_1_data_47),
    .io_rd_small_0_0_data_0(RAMGroup_io_rd_small_0_0_data_0),
    .io_rd_small_0_0_data_1(RAMGroup_io_rd_small_0_0_data_1),
    .io_rd_small_0_0_data_2(RAMGroup_io_rd_small_0_0_data_2),
    .io_rd_small_0_0_data_3(RAMGroup_io_rd_small_0_0_data_3),
    .io_rd_small_0_0_data_4(RAMGroup_io_rd_small_0_0_data_4),
    .io_rd_small_0_0_data_5(RAMGroup_io_rd_small_0_0_data_5),
    .io_rd_small_0_0_data_6(RAMGroup_io_rd_small_0_0_data_6),
    .io_rd_small_0_0_data_7(RAMGroup_io_rd_small_0_0_data_7),
    .io_rd_small_0_1_data_0(RAMGroup_io_rd_small_0_1_data_0),
    .io_rd_small_0_1_data_1(RAMGroup_io_rd_small_0_1_data_1),
    .io_rd_small_0_1_data_2(RAMGroup_io_rd_small_0_1_data_2),
    .io_rd_small_0_1_data_3(RAMGroup_io_rd_small_0_1_data_3),
    .io_rd_small_0_1_data_4(RAMGroup_io_rd_small_0_1_data_4),
    .io_rd_small_0_1_data_5(RAMGroup_io_rd_small_0_1_data_5),
    .io_rd_small_0_1_data_6(RAMGroup_io_rd_small_0_1_data_6),
    .io_rd_small_0_1_data_7(RAMGroup_io_rd_small_0_1_data_7),
    .io_rd_small_0_2_data_0(RAMGroup_io_rd_small_0_2_data_0),
    .io_rd_small_0_2_data_1(RAMGroup_io_rd_small_0_2_data_1),
    .io_rd_small_0_2_data_2(RAMGroup_io_rd_small_0_2_data_2),
    .io_rd_small_0_2_data_3(RAMGroup_io_rd_small_0_2_data_3),
    .io_rd_small_0_2_data_4(RAMGroup_io_rd_small_0_2_data_4),
    .io_rd_small_0_2_data_5(RAMGroup_io_rd_small_0_2_data_5),
    .io_rd_small_0_2_data_6(RAMGroup_io_rd_small_0_2_data_6),
    .io_rd_small_0_2_data_7(RAMGroup_io_rd_small_0_2_data_7),
    .io_rd_small_0_3_data_0(RAMGroup_io_rd_small_0_3_data_0),
    .io_rd_small_0_3_data_1(RAMGroup_io_rd_small_0_3_data_1),
    .io_rd_small_0_3_data_2(RAMGroup_io_rd_small_0_3_data_2),
    .io_rd_small_0_3_data_3(RAMGroup_io_rd_small_0_3_data_3),
    .io_rd_small_0_3_data_4(RAMGroup_io_rd_small_0_3_data_4),
    .io_rd_small_0_3_data_5(RAMGroup_io_rd_small_0_3_data_5),
    .io_rd_small_0_3_data_6(RAMGroup_io_rd_small_0_3_data_6),
    .io_rd_small_0_3_data_7(RAMGroup_io_rd_small_0_3_data_7),
    .io_rd_small_1_0_data_0(RAMGroup_io_rd_small_1_0_data_0),
    .io_rd_small_1_0_data_1(RAMGroup_io_rd_small_1_0_data_1),
    .io_rd_small_1_0_data_2(RAMGroup_io_rd_small_1_0_data_2),
    .io_rd_small_1_0_data_3(RAMGroup_io_rd_small_1_0_data_3),
    .io_rd_small_1_0_data_4(RAMGroup_io_rd_small_1_0_data_4),
    .io_rd_small_1_0_data_5(RAMGroup_io_rd_small_1_0_data_5),
    .io_rd_small_1_0_data_6(RAMGroup_io_rd_small_1_0_data_6),
    .io_rd_small_1_0_data_7(RAMGroup_io_rd_small_1_0_data_7),
    .io_rd_small_1_1_data_0(RAMGroup_io_rd_small_1_1_data_0),
    .io_rd_small_1_1_data_1(RAMGroup_io_rd_small_1_1_data_1),
    .io_rd_small_1_1_data_2(RAMGroup_io_rd_small_1_1_data_2),
    .io_rd_small_1_1_data_3(RAMGroup_io_rd_small_1_1_data_3),
    .io_rd_small_1_1_data_4(RAMGroup_io_rd_small_1_1_data_4),
    .io_rd_small_1_1_data_5(RAMGroup_io_rd_small_1_1_data_5),
    .io_rd_small_1_1_data_6(RAMGroup_io_rd_small_1_1_data_6),
    .io_rd_small_1_1_data_7(RAMGroup_io_rd_small_1_1_data_7),
    .io_rd_small_1_2_data_0(RAMGroup_io_rd_small_1_2_data_0),
    .io_rd_small_1_2_data_1(RAMGroup_io_rd_small_1_2_data_1),
    .io_rd_small_1_2_data_2(RAMGroup_io_rd_small_1_2_data_2),
    .io_rd_small_1_2_data_3(RAMGroup_io_rd_small_1_2_data_3),
    .io_rd_small_1_2_data_4(RAMGroup_io_rd_small_1_2_data_4),
    .io_rd_small_1_2_data_5(RAMGroup_io_rd_small_1_2_data_5),
    .io_rd_small_1_2_data_6(RAMGroup_io_rd_small_1_2_data_6),
    .io_rd_small_1_2_data_7(RAMGroup_io_rd_small_1_2_data_7),
    .io_rd_small_1_3_data_0(RAMGroup_io_rd_small_1_3_data_0),
    .io_rd_small_1_3_data_1(RAMGroup_io_rd_small_1_3_data_1),
    .io_rd_small_1_3_data_2(RAMGroup_io_rd_small_1_3_data_2),
    .io_rd_small_1_3_data_3(RAMGroup_io_rd_small_1_3_data_3),
    .io_rd_small_1_3_data_4(RAMGroup_io_rd_small_1_3_data_4),
    .io_rd_small_1_3_data_5(RAMGroup_io_rd_small_1_3_data_5),
    .io_rd_small_1_3_data_6(RAMGroup_io_rd_small_1_3_data_6),
    .io_rd_small_1_3_data_7(RAMGroup_io_rd_small_1_3_data_7)
  );
  assign io_complete = 1'h0; // @[top.scala 30:17]
  assign GraphReader_clock = clock;
  assign GraphReader_reset = reset;
  assign GraphReader_io_valid_in = _T ? 1'h0 : _T_1; // @[Conditional.scala 40:58 top.scala 33:22]
  assign GraphReader_io_flag_job = 3'h0 == state; // @[Conditional.scala 37:30]
  assign GraphReader_io_job_big_bank_id = 3'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_big_cnt_x_end = _T ? 10'h3 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_big_cnt_y_end = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_big_cnt_ic_end = _T ? 10'h3 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_big_cnt_loop_end = _T ? 10'h1f : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_big_begin_loop = _T ? 10'h10 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_small_0_max_addr = _T ? 10'h1c1 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_small_0_cnt_y_end = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_small_0_cnt_ic_end = _T ? 10'h3 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_small_0_cnt_loop_end = _T ? 10'h1f : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_small_0_begin_loop = _T ? 10'h10 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_io_job_small_0_cnt_invalid_end = _T ? 10'h100 : 10'h0; // @[Conditional.scala 40:58 para.scala 39:21 top.scala 34:17]
  assign GraphReader_1_clock = clock;
  assign GraphReader_1_reset = reset;
  assign GraphReader_1_io_valid_in = _T ? 1'h0 : _T_1; // @[Conditional.scala 40:58 top.scala 33:22]
  assign GraphReader_1_io_flag_job = 3'h0 == state; // @[Conditional.scala 37:30]
  assign GraphReader_1_io_job_big_bank_id = _T ? 3'h1 : 3'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_big_cnt_x_end = _T ? 10'h3 : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_big_cnt_y_end = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_big_cnt_ic_end = _T ? 10'h3 : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_big_cnt_loop_end = _T ? 10'h1f : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_big_begin_loop = 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_small_0_max_addr = _T ? 10'h1c1 : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_small_0_cnt_y_end = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_small_0_cnt_ic_end = _T ? 10'h3 : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_small_0_cnt_loop_end = _T ? 10'h1f : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_small_0_begin_loop = 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign GraphReader_1_io_job_small_0_cnt_invalid_end = _T ? 10'h100 : 10'h0; // @[Conditional.scala 40:58 para.scala 58:21 top.scala 41:17]
  assign PackReadData_clock = clock;
  assign PackReadData_reset = reset;
  assign PackReadData_io_valid_in = RAMGroup_io_rd_valid_out; // @[top.scala 51:24]
  assign PackReadData_io_flag_job = 3'h0 == state; // @[Conditional.scala 37:30]
  assign PackReadData_io_job_cnt_x_end = _T ? 10'h3 : 10'h0; // @[Conditional.scala 40:58 para.scala 80:16 top.scala 53:19]
  assign PackReadData_io_job_cnt_y_end = _T ? 10'h3 : 10'h0; // @[Conditional.scala 40:58 para.scala 80:16 top.scala 53:19]
  assign PackReadData_io_job_in_chan = _T ? 10'h3f : 10'h0; // @[Conditional.scala 40:58 para.scala 80:16 top.scala 53:19]
  assign PackReadData_io_from_big_0_data_0 = RAMGroup_io_rd_big_0_data_0; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_1 = RAMGroup_io_rd_big_0_data_1; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_2 = RAMGroup_io_rd_big_0_data_2; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_3 = RAMGroup_io_rd_big_0_data_3; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_4 = RAMGroup_io_rd_big_0_data_4; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_5 = RAMGroup_io_rd_big_0_data_5; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_6 = RAMGroup_io_rd_big_0_data_6; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_7 = RAMGroup_io_rd_big_0_data_7; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_8 = RAMGroup_io_rd_big_0_data_8; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_9 = RAMGroup_io_rd_big_0_data_9; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_10 = RAMGroup_io_rd_big_0_data_10; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_11 = RAMGroup_io_rd_big_0_data_11; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_12 = RAMGroup_io_rd_big_0_data_12; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_13 = RAMGroup_io_rd_big_0_data_13; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_14 = RAMGroup_io_rd_big_0_data_14; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_15 = RAMGroup_io_rd_big_0_data_15; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_16 = RAMGroup_io_rd_big_0_data_16; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_17 = RAMGroup_io_rd_big_0_data_17; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_18 = RAMGroup_io_rd_big_0_data_18; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_19 = RAMGroup_io_rd_big_0_data_19; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_20 = RAMGroup_io_rd_big_0_data_20; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_21 = RAMGroup_io_rd_big_0_data_21; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_22 = RAMGroup_io_rd_big_0_data_22; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_23 = RAMGroup_io_rd_big_0_data_23; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_24 = RAMGroup_io_rd_big_0_data_24; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_25 = RAMGroup_io_rd_big_0_data_25; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_26 = RAMGroup_io_rd_big_0_data_26; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_27 = RAMGroup_io_rd_big_0_data_27; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_28 = RAMGroup_io_rd_big_0_data_28; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_29 = RAMGroup_io_rd_big_0_data_29; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_30 = RAMGroup_io_rd_big_0_data_30; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_31 = RAMGroup_io_rd_big_0_data_31; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_32 = RAMGroup_io_rd_big_0_data_32; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_33 = RAMGroup_io_rd_big_0_data_33; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_34 = RAMGroup_io_rd_big_0_data_34; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_35 = RAMGroup_io_rd_big_0_data_35; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_36 = RAMGroup_io_rd_big_0_data_36; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_37 = RAMGroup_io_rd_big_0_data_37; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_38 = RAMGroup_io_rd_big_0_data_38; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_39 = RAMGroup_io_rd_big_0_data_39; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_40 = RAMGroup_io_rd_big_0_data_40; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_41 = RAMGroup_io_rd_big_0_data_41; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_42 = RAMGroup_io_rd_big_0_data_42; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_43 = RAMGroup_io_rd_big_0_data_43; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_44 = RAMGroup_io_rd_big_0_data_44; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_45 = RAMGroup_io_rd_big_0_data_45; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_46 = RAMGroup_io_rd_big_0_data_46; // @[top.scala 54:24]
  assign PackReadData_io_from_big_0_data_47 = RAMGroup_io_rd_big_0_data_47; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_0 = RAMGroup_io_rd_big_1_data_0; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_1 = RAMGroup_io_rd_big_1_data_1; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_2 = RAMGroup_io_rd_big_1_data_2; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_3 = RAMGroup_io_rd_big_1_data_3; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_4 = RAMGroup_io_rd_big_1_data_4; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_5 = RAMGroup_io_rd_big_1_data_5; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_6 = RAMGroup_io_rd_big_1_data_6; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_7 = RAMGroup_io_rd_big_1_data_7; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_8 = RAMGroup_io_rd_big_1_data_8; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_9 = RAMGroup_io_rd_big_1_data_9; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_10 = RAMGroup_io_rd_big_1_data_10; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_11 = RAMGroup_io_rd_big_1_data_11; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_12 = RAMGroup_io_rd_big_1_data_12; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_13 = RAMGroup_io_rd_big_1_data_13; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_14 = RAMGroup_io_rd_big_1_data_14; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_15 = RAMGroup_io_rd_big_1_data_15; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_16 = RAMGroup_io_rd_big_1_data_16; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_17 = RAMGroup_io_rd_big_1_data_17; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_18 = RAMGroup_io_rd_big_1_data_18; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_19 = RAMGroup_io_rd_big_1_data_19; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_20 = RAMGroup_io_rd_big_1_data_20; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_21 = RAMGroup_io_rd_big_1_data_21; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_22 = RAMGroup_io_rd_big_1_data_22; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_23 = RAMGroup_io_rd_big_1_data_23; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_24 = RAMGroup_io_rd_big_1_data_24; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_25 = RAMGroup_io_rd_big_1_data_25; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_26 = RAMGroup_io_rd_big_1_data_26; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_27 = RAMGroup_io_rd_big_1_data_27; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_28 = RAMGroup_io_rd_big_1_data_28; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_29 = RAMGroup_io_rd_big_1_data_29; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_30 = RAMGroup_io_rd_big_1_data_30; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_31 = RAMGroup_io_rd_big_1_data_31; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_32 = RAMGroup_io_rd_big_1_data_32; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_33 = RAMGroup_io_rd_big_1_data_33; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_34 = RAMGroup_io_rd_big_1_data_34; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_35 = RAMGroup_io_rd_big_1_data_35; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_36 = RAMGroup_io_rd_big_1_data_36; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_37 = RAMGroup_io_rd_big_1_data_37; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_38 = RAMGroup_io_rd_big_1_data_38; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_39 = RAMGroup_io_rd_big_1_data_39; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_40 = RAMGroup_io_rd_big_1_data_40; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_41 = RAMGroup_io_rd_big_1_data_41; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_42 = RAMGroup_io_rd_big_1_data_42; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_43 = RAMGroup_io_rd_big_1_data_43; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_44 = RAMGroup_io_rd_big_1_data_44; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_45 = RAMGroup_io_rd_big_1_data_45; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_46 = RAMGroup_io_rd_big_1_data_46; // @[top.scala 54:24]
  assign PackReadData_io_from_big_1_data_47 = RAMGroup_io_rd_big_1_data_47; // @[top.scala 54:24]
  assign PackReadData_io_from_small_0_0_data_0 = RAMGroup_io_rd_small_0_0_data_0; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_0_data_1 = RAMGroup_io_rd_small_0_0_data_1; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_0_data_2 = RAMGroup_io_rd_small_0_0_data_2; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_0_data_3 = RAMGroup_io_rd_small_0_0_data_3; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_0_data_4 = RAMGroup_io_rd_small_0_0_data_4; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_0_data_5 = RAMGroup_io_rd_small_0_0_data_5; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_0_data_6 = RAMGroup_io_rd_small_0_0_data_6; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_0_data_7 = RAMGroup_io_rd_small_0_0_data_7; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_1_data_0 = RAMGroup_io_rd_small_0_1_data_0; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_1_data_1 = RAMGroup_io_rd_small_0_1_data_1; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_1_data_2 = RAMGroup_io_rd_small_0_1_data_2; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_1_data_3 = RAMGroup_io_rd_small_0_1_data_3; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_1_data_4 = RAMGroup_io_rd_small_0_1_data_4; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_1_data_5 = RAMGroup_io_rd_small_0_1_data_5; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_1_data_6 = RAMGroup_io_rd_small_0_1_data_6; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_1_data_7 = RAMGroup_io_rd_small_0_1_data_7; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_2_data_0 = RAMGroup_io_rd_small_0_2_data_0; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_2_data_1 = RAMGroup_io_rd_small_0_2_data_1; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_2_data_2 = RAMGroup_io_rd_small_0_2_data_2; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_2_data_3 = RAMGroup_io_rd_small_0_2_data_3; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_2_data_4 = RAMGroup_io_rd_small_0_2_data_4; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_2_data_5 = RAMGroup_io_rd_small_0_2_data_5; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_2_data_6 = RAMGroup_io_rd_small_0_2_data_6; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_2_data_7 = RAMGroup_io_rd_small_0_2_data_7; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_3_data_0 = RAMGroup_io_rd_small_0_3_data_0; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_3_data_1 = RAMGroup_io_rd_small_0_3_data_1; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_3_data_2 = RAMGroup_io_rd_small_0_3_data_2; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_3_data_3 = RAMGroup_io_rd_small_0_3_data_3; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_3_data_4 = RAMGroup_io_rd_small_0_3_data_4; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_3_data_5 = RAMGroup_io_rd_small_0_3_data_5; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_3_data_6 = RAMGroup_io_rd_small_0_3_data_6; // @[top.scala 55:26]
  assign PackReadData_io_from_small_0_3_data_7 = RAMGroup_io_rd_small_0_3_data_7; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_0_data_0 = RAMGroup_io_rd_small_1_0_data_0; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_0_data_1 = RAMGroup_io_rd_small_1_0_data_1; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_0_data_2 = RAMGroup_io_rd_small_1_0_data_2; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_0_data_3 = RAMGroup_io_rd_small_1_0_data_3; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_0_data_4 = RAMGroup_io_rd_small_1_0_data_4; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_0_data_5 = RAMGroup_io_rd_small_1_0_data_5; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_0_data_6 = RAMGroup_io_rd_small_1_0_data_6; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_0_data_7 = RAMGroup_io_rd_small_1_0_data_7; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_1_data_0 = RAMGroup_io_rd_small_1_1_data_0; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_1_data_1 = RAMGroup_io_rd_small_1_1_data_1; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_1_data_2 = RAMGroup_io_rd_small_1_1_data_2; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_1_data_3 = RAMGroup_io_rd_small_1_1_data_3; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_1_data_4 = RAMGroup_io_rd_small_1_1_data_4; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_1_data_5 = RAMGroup_io_rd_small_1_1_data_5; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_1_data_6 = RAMGroup_io_rd_small_1_1_data_6; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_1_data_7 = RAMGroup_io_rd_small_1_1_data_7; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_2_data_0 = RAMGroup_io_rd_small_1_2_data_0; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_2_data_1 = RAMGroup_io_rd_small_1_2_data_1; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_2_data_2 = RAMGroup_io_rd_small_1_2_data_2; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_2_data_3 = RAMGroup_io_rd_small_1_2_data_3; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_2_data_4 = RAMGroup_io_rd_small_1_2_data_4; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_2_data_5 = RAMGroup_io_rd_small_1_2_data_5; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_2_data_6 = RAMGroup_io_rd_small_1_2_data_6; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_2_data_7 = RAMGroup_io_rd_small_1_2_data_7; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_3_data_0 = RAMGroup_io_rd_small_1_3_data_0; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_3_data_1 = RAMGroup_io_rd_small_1_3_data_1; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_3_data_2 = RAMGroup_io_rd_small_1_3_data_2; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_3_data_3 = RAMGroup_io_rd_small_1_3_data_3; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_3_data_4 = RAMGroup_io_rd_small_1_3_data_4; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_3_data_5 = RAMGroup_io_rd_small_1_3_data_5; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_3_data_6 = RAMGroup_io_rd_small_1_3_data_6; // @[top.scala 55:26]
  assign PackReadData_io_from_small_1_3_data_7 = RAMGroup_io_rd_small_1_3_data_7; // @[top.scala 55:26]
  assign ReadSwitch_clock = clock;
  assign ReadSwitch_reset = reset;
  assign ReadSwitch_io_flag_job = 3'h0 == state; // @[Conditional.scala 37:30]
  assign ReadSwitch_io_job = _T ? 2'h1 : 2'h0; // @[Conditional.scala 40:58 para.scala 86:16 top.scala 58:21]
  assign ReadSwitch_io_valid_in = PackReadData_io_valid_out; // @[top.scala 59:26]
  assign ReadSwitch_io_from_mat_0 = PackReadData_io_output_mat_0; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_1 = PackReadData_io_output_mat_1; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_2 = PackReadData_io_output_mat_2; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_3 = PackReadData_io_output_mat_3; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_4 = PackReadData_io_output_mat_4; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_5 = PackReadData_io_output_mat_5; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_6 = PackReadData_io_output_mat_6; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_7 = PackReadData_io_output_mat_7; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_8 = PackReadData_io_output_mat_8; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_9 = PackReadData_io_output_mat_9; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_10 = PackReadData_io_output_mat_10; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_11 = PackReadData_io_output_mat_11; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_12 = PackReadData_io_output_mat_12; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_13 = PackReadData_io_output_mat_13; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_14 = PackReadData_io_output_mat_14; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_15 = PackReadData_io_output_mat_15; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_16 = PackReadData_io_output_mat_16; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_17 = PackReadData_io_output_mat_17; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_18 = PackReadData_io_output_mat_18; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_19 = PackReadData_io_output_mat_19; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_20 = PackReadData_io_output_mat_20; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_21 = PackReadData_io_output_mat_21; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_22 = PackReadData_io_output_mat_22; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_23 = PackReadData_io_output_mat_23; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_24 = PackReadData_io_output_mat_24; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_25 = PackReadData_io_output_mat_25; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_26 = PackReadData_io_output_mat_26; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_27 = PackReadData_io_output_mat_27; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_28 = PackReadData_io_output_mat_28; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_29 = PackReadData_io_output_mat_29; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_30 = PackReadData_io_output_mat_30; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_31 = PackReadData_io_output_mat_31; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_32 = PackReadData_io_output_mat_32; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_33 = PackReadData_io_output_mat_33; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_34 = PackReadData_io_output_mat_34; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_35 = PackReadData_io_output_mat_35; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_36 = PackReadData_io_output_mat_36; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_37 = PackReadData_io_output_mat_37; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_38 = PackReadData_io_output_mat_38; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_39 = PackReadData_io_output_mat_39; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_40 = PackReadData_io_output_mat_40; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_41 = PackReadData_io_output_mat_41; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_42 = PackReadData_io_output_mat_42; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_43 = PackReadData_io_output_mat_43; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_44 = PackReadData_io_output_mat_44; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_45 = PackReadData_io_output_mat_45; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_46 = PackReadData_io_output_mat_46; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_47 = PackReadData_io_output_mat_47; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_48 = PackReadData_io_output_mat_48; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_49 = PackReadData_io_output_mat_49; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_50 = PackReadData_io_output_mat_50; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_51 = PackReadData_io_output_mat_51; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_52 = PackReadData_io_output_mat_52; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_53 = PackReadData_io_output_mat_53; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_54 = PackReadData_io_output_mat_54; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_55 = PackReadData_io_output_mat_55; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_56 = PackReadData_io_output_mat_56; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_57 = PackReadData_io_output_mat_57; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_58 = PackReadData_io_output_mat_58; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_59 = PackReadData_io_output_mat_59; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_60 = PackReadData_io_output_mat_60; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_61 = PackReadData_io_output_mat_61; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_62 = PackReadData_io_output_mat_62; // @[top.scala 60:22]
  assign ReadSwitch_io_from_mat_63 = PackReadData_io_output_mat_63; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_0 = PackReadData_io_output_up_0; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_1 = PackReadData_io_output_up_1; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_2 = PackReadData_io_output_up_2; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_3 = PackReadData_io_output_up_3; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_4 = PackReadData_io_output_up_4; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_5 = PackReadData_io_output_up_5; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_6 = PackReadData_io_output_up_6; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_7 = PackReadData_io_output_up_7; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_8 = PackReadData_io_output_up_8; // @[top.scala 60:22]
  assign ReadSwitch_io_from_up_9 = PackReadData_io_output_up_9; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_0 = PackReadData_io_output_down_0; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_1 = PackReadData_io_output_down_1; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_2 = PackReadData_io_output_down_2; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_3 = PackReadData_io_output_down_3; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_4 = PackReadData_io_output_down_4; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_5 = PackReadData_io_output_down_5; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_6 = PackReadData_io_output_down_6; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_7 = PackReadData_io_output_down_7; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_8 = PackReadData_io_output_down_8; // @[top.scala 60:22]
  assign ReadSwitch_io_from_down_9 = PackReadData_io_output_down_9; // @[top.scala 60:22]
  assign ReadSwitch_io_from_left_0 = PackReadData_io_output_left_0; // @[top.scala 60:22]
  assign ReadSwitch_io_from_left_1 = PackReadData_io_output_left_1; // @[top.scala 60:22]
  assign ReadSwitch_io_from_left_2 = PackReadData_io_output_left_2; // @[top.scala 60:22]
  assign ReadSwitch_io_from_left_3 = PackReadData_io_output_left_3; // @[top.scala 60:22]
  assign ReadSwitch_io_from_left_4 = PackReadData_io_output_left_4; // @[top.scala 60:22]
  assign ReadSwitch_io_from_left_5 = PackReadData_io_output_left_5; // @[top.scala 60:22]
  assign ReadSwitch_io_from_left_6 = PackReadData_io_output_left_6; // @[top.scala 60:22]
  assign ReadSwitch_io_from_left_7 = PackReadData_io_output_left_7; // @[top.scala 60:22]
  assign ReadSwitch_io_from_right_0 = PackReadData_io_output_right_0; // @[top.scala 60:22]
  assign ReadSwitch_io_from_right_1 = PackReadData_io_output_right_1; // @[top.scala 60:22]
  assign ReadSwitch_io_from_right_2 = PackReadData_io_output_right_2; // @[top.scala 60:22]
  assign ReadSwitch_io_from_right_3 = PackReadData_io_output_right_3; // @[top.scala 60:22]
  assign ReadSwitch_io_from_right_4 = PackReadData_io_output_right_4; // @[top.scala 60:22]
  assign ReadSwitch_io_from_right_5 = PackReadData_io_output_right_5; // @[top.scala 60:22]
  assign ReadSwitch_io_from_right_6 = PackReadData_io_output_right_6; // @[top.scala 60:22]
  assign ReadSwitch_io_from_right_7 = PackReadData_io_output_right_7; // @[top.scala 60:22]
  assign ReadSwitch_io_from_weight_0 = ROMWeight_io_out_0; // @[top.scala 61:29]
  assign ReadSwitch_io_from_weight_1 = ROMWeight_io_out_1; // @[top.scala 61:29]
  assign ReadSwitch_io_from_weight_2 = ROMWeight_io_out_2; // @[top.scala 61:29]
  assign ReadSwitch_io_from_weight_3 = ROMWeight_io_out_3; // @[top.scala 61:29]
  assign ReadSwitch_io_from_weight_4 = ROMWeight_io_out_4; // @[top.scala 61:29]
  assign ReadSwitch_io_from_weight_5 = ROMWeight_io_out_5; // @[top.scala 61:29]
  assign ReadSwitch_io_from_weight_6 = ROMWeight_io_out_6; // @[top.scala 61:29]
  assign ReadSwitch_io_from_weight_7 = ROMWeight_io_out_7; // @[top.scala 61:29]
  assign ReadSwitch_io_from_weight_8 = ROMWeight_io_out_8; // @[top.scala 61:29]
  assign WeightReader_clock = clock;
  assign WeightReader_reset = reset;
  assign WeightReader_io_valid_in = _T ? 1'h0 : _T_1; // @[Conditional.scala 40:58 top.scala 33:22]
  assign WeightReader_io_flag_job = 3'h0 == state; // @[Conditional.scala 37:30]
  assign WeightReader_io_addr_end = {{8'd0}, _GEN_148}; // @[Conditional.scala 40:58 para.scala 74:21 top.scala 45:26]
  assign Calc8x8_clock = clock;
  assign Calc8x8_reset = reset;
  assign Calc8x8_io_input_mat_0 = ReadSwitch_io_to_calc8x8_mat_0; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_1 = ReadSwitch_io_to_calc8x8_mat_1; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_2 = ReadSwitch_io_to_calc8x8_mat_2; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_3 = ReadSwitch_io_to_calc8x8_mat_3; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_4 = ReadSwitch_io_to_calc8x8_mat_4; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_5 = ReadSwitch_io_to_calc8x8_mat_5; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_6 = ReadSwitch_io_to_calc8x8_mat_6; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_7 = ReadSwitch_io_to_calc8x8_mat_7; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_8 = ReadSwitch_io_to_calc8x8_mat_8; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_9 = ReadSwitch_io_to_calc8x8_mat_9; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_10 = ReadSwitch_io_to_calc8x8_mat_10; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_11 = ReadSwitch_io_to_calc8x8_mat_11; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_12 = ReadSwitch_io_to_calc8x8_mat_12; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_13 = ReadSwitch_io_to_calc8x8_mat_13; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_14 = ReadSwitch_io_to_calc8x8_mat_14; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_15 = ReadSwitch_io_to_calc8x8_mat_15; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_16 = ReadSwitch_io_to_calc8x8_mat_16; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_17 = ReadSwitch_io_to_calc8x8_mat_17; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_18 = ReadSwitch_io_to_calc8x8_mat_18; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_19 = ReadSwitch_io_to_calc8x8_mat_19; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_20 = ReadSwitch_io_to_calc8x8_mat_20; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_21 = ReadSwitch_io_to_calc8x8_mat_21; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_22 = ReadSwitch_io_to_calc8x8_mat_22; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_23 = ReadSwitch_io_to_calc8x8_mat_23; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_24 = ReadSwitch_io_to_calc8x8_mat_24; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_25 = ReadSwitch_io_to_calc8x8_mat_25; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_26 = ReadSwitch_io_to_calc8x8_mat_26; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_27 = ReadSwitch_io_to_calc8x8_mat_27; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_28 = ReadSwitch_io_to_calc8x8_mat_28; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_29 = ReadSwitch_io_to_calc8x8_mat_29; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_30 = ReadSwitch_io_to_calc8x8_mat_30; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_31 = ReadSwitch_io_to_calc8x8_mat_31; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_32 = ReadSwitch_io_to_calc8x8_mat_32; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_33 = ReadSwitch_io_to_calc8x8_mat_33; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_34 = ReadSwitch_io_to_calc8x8_mat_34; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_35 = ReadSwitch_io_to_calc8x8_mat_35; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_36 = ReadSwitch_io_to_calc8x8_mat_36; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_37 = ReadSwitch_io_to_calc8x8_mat_37; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_38 = ReadSwitch_io_to_calc8x8_mat_38; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_39 = ReadSwitch_io_to_calc8x8_mat_39; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_40 = ReadSwitch_io_to_calc8x8_mat_40; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_41 = ReadSwitch_io_to_calc8x8_mat_41; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_42 = ReadSwitch_io_to_calc8x8_mat_42; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_43 = ReadSwitch_io_to_calc8x8_mat_43; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_44 = ReadSwitch_io_to_calc8x8_mat_44; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_45 = ReadSwitch_io_to_calc8x8_mat_45; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_46 = ReadSwitch_io_to_calc8x8_mat_46; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_47 = ReadSwitch_io_to_calc8x8_mat_47; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_48 = ReadSwitch_io_to_calc8x8_mat_48; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_49 = ReadSwitch_io_to_calc8x8_mat_49; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_50 = ReadSwitch_io_to_calc8x8_mat_50; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_51 = ReadSwitch_io_to_calc8x8_mat_51; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_52 = ReadSwitch_io_to_calc8x8_mat_52; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_53 = ReadSwitch_io_to_calc8x8_mat_53; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_54 = ReadSwitch_io_to_calc8x8_mat_54; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_55 = ReadSwitch_io_to_calc8x8_mat_55; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_56 = ReadSwitch_io_to_calc8x8_mat_56; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_57 = ReadSwitch_io_to_calc8x8_mat_57; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_58 = ReadSwitch_io_to_calc8x8_mat_58; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_59 = ReadSwitch_io_to_calc8x8_mat_59; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_60 = ReadSwitch_io_to_calc8x8_mat_60; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_61 = ReadSwitch_io_to_calc8x8_mat_61; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_62 = ReadSwitch_io_to_calc8x8_mat_62; // @[top.scala 63:19]
  assign Calc8x8_io_input_mat_63 = ReadSwitch_io_to_calc8x8_mat_63; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_0 = ReadSwitch_io_to_calc8x8_up_0; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_1 = ReadSwitch_io_to_calc8x8_up_1; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_2 = ReadSwitch_io_to_calc8x8_up_2; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_3 = ReadSwitch_io_to_calc8x8_up_3; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_4 = ReadSwitch_io_to_calc8x8_up_4; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_5 = ReadSwitch_io_to_calc8x8_up_5; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_6 = ReadSwitch_io_to_calc8x8_up_6; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_7 = ReadSwitch_io_to_calc8x8_up_7; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_8 = ReadSwitch_io_to_calc8x8_up_8; // @[top.scala 63:19]
  assign Calc8x8_io_input_up_9 = ReadSwitch_io_to_calc8x8_up_9; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_0 = ReadSwitch_io_to_calc8x8_down_0; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_1 = ReadSwitch_io_to_calc8x8_down_1; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_2 = ReadSwitch_io_to_calc8x8_down_2; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_3 = ReadSwitch_io_to_calc8x8_down_3; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_4 = ReadSwitch_io_to_calc8x8_down_4; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_5 = ReadSwitch_io_to_calc8x8_down_5; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_6 = ReadSwitch_io_to_calc8x8_down_6; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_7 = ReadSwitch_io_to_calc8x8_down_7; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_8 = ReadSwitch_io_to_calc8x8_down_8; // @[top.scala 63:19]
  assign Calc8x8_io_input_down_9 = ReadSwitch_io_to_calc8x8_down_9; // @[top.scala 63:19]
  assign Calc8x8_io_input_left_0 = ReadSwitch_io_to_calc8x8_left_0; // @[top.scala 63:19]
  assign Calc8x8_io_input_left_1 = ReadSwitch_io_to_calc8x8_left_1; // @[top.scala 63:19]
  assign Calc8x8_io_input_left_2 = ReadSwitch_io_to_calc8x8_left_2; // @[top.scala 63:19]
  assign Calc8x8_io_input_left_3 = ReadSwitch_io_to_calc8x8_left_3; // @[top.scala 63:19]
  assign Calc8x8_io_input_left_4 = ReadSwitch_io_to_calc8x8_left_4; // @[top.scala 63:19]
  assign Calc8x8_io_input_left_5 = ReadSwitch_io_to_calc8x8_left_5; // @[top.scala 63:19]
  assign Calc8x8_io_input_left_6 = ReadSwitch_io_to_calc8x8_left_6; // @[top.scala 63:19]
  assign Calc8x8_io_input_left_7 = ReadSwitch_io_to_calc8x8_left_7; // @[top.scala 63:19]
  assign Calc8x8_io_input_right_0 = ReadSwitch_io_to_calc8x8_right_0; // @[top.scala 63:19]
  assign Calc8x8_io_input_right_1 = ReadSwitch_io_to_calc8x8_right_1; // @[top.scala 63:19]
  assign Calc8x8_io_input_right_2 = ReadSwitch_io_to_calc8x8_right_2; // @[top.scala 63:19]
  assign Calc8x8_io_input_right_3 = ReadSwitch_io_to_calc8x8_right_3; // @[top.scala 63:19]
  assign Calc8x8_io_input_right_4 = ReadSwitch_io_to_calc8x8_right_4; // @[top.scala 63:19]
  assign Calc8x8_io_input_right_5 = ReadSwitch_io_to_calc8x8_right_5; // @[top.scala 63:19]
  assign Calc8x8_io_input_right_6 = ReadSwitch_io_to_calc8x8_right_6; // @[top.scala 63:19]
  assign Calc8x8_io_input_right_7 = ReadSwitch_io_to_calc8x8_right_7; // @[top.scala 63:19]
  assign Calc8x8_io_flag = _T ? 2'h2 : _GEN_7; // @[Conditional.scala 40:58 top.scala 147:26]
  assign Calc8x8_io_weight_0_real_0 = ReadSwitch_io_to_weight_0_real_0; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_1 = ReadSwitch_io_to_weight_0_real_1; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_2 = ReadSwitch_io_to_weight_0_real_2; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_3 = ReadSwitch_io_to_weight_0_real_3; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_4 = ReadSwitch_io_to_weight_0_real_4; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_5 = ReadSwitch_io_to_weight_0_real_5; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_6 = ReadSwitch_io_to_weight_0_real_6; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_7 = ReadSwitch_io_to_weight_0_real_7; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_8 = ReadSwitch_io_to_weight_0_real_8; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_9 = ReadSwitch_io_to_weight_0_real_9; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_10 = ReadSwitch_io_to_weight_0_real_10; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_11 = ReadSwitch_io_to_weight_0_real_11; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_12 = ReadSwitch_io_to_weight_0_real_12; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_13 = ReadSwitch_io_to_weight_0_real_13; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_14 = ReadSwitch_io_to_weight_0_real_14; // @[top.scala 65:20]
  assign Calc8x8_io_weight_0_real_15 = ReadSwitch_io_to_weight_0_real_15; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_0 = ReadSwitch_io_to_weight_1_real_0; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_1 = ReadSwitch_io_to_weight_1_real_1; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_2 = ReadSwitch_io_to_weight_1_real_2; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_3 = ReadSwitch_io_to_weight_1_real_3; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_4 = ReadSwitch_io_to_weight_1_real_4; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_5 = ReadSwitch_io_to_weight_1_real_5; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_6 = ReadSwitch_io_to_weight_1_real_6; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_7 = ReadSwitch_io_to_weight_1_real_7; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_8 = ReadSwitch_io_to_weight_1_real_8; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_9 = ReadSwitch_io_to_weight_1_real_9; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_10 = ReadSwitch_io_to_weight_1_real_10; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_11 = ReadSwitch_io_to_weight_1_real_11; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_12 = ReadSwitch_io_to_weight_1_real_12; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_13 = ReadSwitch_io_to_weight_1_real_13; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_14 = ReadSwitch_io_to_weight_1_real_14; // @[top.scala 65:20]
  assign Calc8x8_io_weight_1_real_15 = ReadSwitch_io_to_weight_1_real_15; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_0 = ReadSwitch_io_to_weight_2_real_0; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_1 = ReadSwitch_io_to_weight_2_real_1; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_2 = ReadSwitch_io_to_weight_2_real_2; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_3 = ReadSwitch_io_to_weight_2_real_3; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_4 = ReadSwitch_io_to_weight_2_real_4; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_5 = ReadSwitch_io_to_weight_2_real_5; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_6 = ReadSwitch_io_to_weight_2_real_6; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_7 = ReadSwitch_io_to_weight_2_real_7; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_8 = ReadSwitch_io_to_weight_2_real_8; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_9 = ReadSwitch_io_to_weight_2_real_9; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_10 = ReadSwitch_io_to_weight_2_real_10; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_11 = ReadSwitch_io_to_weight_2_real_11; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_12 = ReadSwitch_io_to_weight_2_real_12; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_13 = ReadSwitch_io_to_weight_2_real_13; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_14 = ReadSwitch_io_to_weight_2_real_14; // @[top.scala 65:20]
  assign Calc8x8_io_weight_2_real_15 = ReadSwitch_io_to_weight_2_real_15; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_0 = ReadSwitch_io_to_weight_3_real_0; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_1 = ReadSwitch_io_to_weight_3_real_1; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_2 = ReadSwitch_io_to_weight_3_real_2; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_3 = ReadSwitch_io_to_weight_3_real_3; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_4 = ReadSwitch_io_to_weight_3_real_4; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_5 = ReadSwitch_io_to_weight_3_real_5; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_6 = ReadSwitch_io_to_weight_3_real_6; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_7 = ReadSwitch_io_to_weight_3_real_7; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_8 = ReadSwitch_io_to_weight_3_real_8; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_9 = ReadSwitch_io_to_weight_3_real_9; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_10 = ReadSwitch_io_to_weight_3_real_10; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_11 = ReadSwitch_io_to_weight_3_real_11; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_12 = ReadSwitch_io_to_weight_3_real_12; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_13 = ReadSwitch_io_to_weight_3_real_13; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_14 = ReadSwitch_io_to_weight_3_real_14; // @[top.scala 65:20]
  assign Calc8x8_io_weight_3_real_15 = ReadSwitch_io_to_weight_3_real_15; // @[top.scala 65:20]
  assign Calc8x8_io_valid_in = ReadSwitch_io_valid_out_calc8x8; // @[top.scala 66:22]
  assign Accumu_clock = clock;
  assign Accumu_reset = reset;
  assign Accumu_io_valid_in = Calc8x8_io_valid_out; // @[top.scala 70:19]
  assign Accumu_io_flag_job = 3'h0 == state; // @[Conditional.scala 37:30]
  assign Accumu_io_in_from_calc8x8_mat_0 = Calc8x8_io_output_mat_0; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_1 = Calc8x8_io_output_mat_1; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_2 = Calc8x8_io_output_mat_2; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_3 = Calc8x8_io_output_mat_3; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_4 = Calc8x8_io_output_mat_4; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_5 = Calc8x8_io_output_mat_5; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_6 = Calc8x8_io_output_mat_6; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_7 = Calc8x8_io_output_mat_7; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_8 = Calc8x8_io_output_mat_8; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_9 = Calc8x8_io_output_mat_9; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_10 = Calc8x8_io_output_mat_10; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_11 = Calc8x8_io_output_mat_11; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_12 = Calc8x8_io_output_mat_12; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_13 = Calc8x8_io_output_mat_13; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_14 = Calc8x8_io_output_mat_14; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_15 = Calc8x8_io_output_mat_15; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_16 = Calc8x8_io_output_mat_16; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_17 = Calc8x8_io_output_mat_17; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_18 = Calc8x8_io_output_mat_18; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_19 = Calc8x8_io_output_mat_19; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_20 = Calc8x8_io_output_mat_20; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_21 = Calc8x8_io_output_mat_21; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_22 = Calc8x8_io_output_mat_22; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_23 = Calc8x8_io_output_mat_23; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_24 = Calc8x8_io_output_mat_24; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_25 = Calc8x8_io_output_mat_25; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_26 = Calc8x8_io_output_mat_26; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_27 = Calc8x8_io_output_mat_27; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_28 = Calc8x8_io_output_mat_28; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_29 = Calc8x8_io_output_mat_29; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_30 = Calc8x8_io_output_mat_30; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_31 = Calc8x8_io_output_mat_31; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_32 = Calc8x8_io_output_mat_32; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_33 = Calc8x8_io_output_mat_33; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_34 = Calc8x8_io_output_mat_34; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_35 = Calc8x8_io_output_mat_35; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_36 = Calc8x8_io_output_mat_36; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_37 = Calc8x8_io_output_mat_37; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_38 = Calc8x8_io_output_mat_38; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_39 = Calc8x8_io_output_mat_39; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_40 = Calc8x8_io_output_mat_40; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_41 = Calc8x8_io_output_mat_41; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_42 = Calc8x8_io_output_mat_42; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_43 = Calc8x8_io_output_mat_43; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_44 = Calc8x8_io_output_mat_44; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_45 = Calc8x8_io_output_mat_45; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_46 = Calc8x8_io_output_mat_46; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_47 = Calc8x8_io_output_mat_47; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_48 = Calc8x8_io_output_mat_48; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_49 = Calc8x8_io_output_mat_49; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_50 = Calc8x8_io_output_mat_50; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_51 = Calc8x8_io_output_mat_51; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_52 = Calc8x8_io_output_mat_52; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_53 = Calc8x8_io_output_mat_53; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_54 = Calc8x8_io_output_mat_54; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_55 = Calc8x8_io_output_mat_55; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_56 = Calc8x8_io_output_mat_56; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_57 = Calc8x8_io_output_mat_57; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_58 = Calc8x8_io_output_mat_58; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_59 = Calc8x8_io_output_mat_59; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_60 = Calc8x8_io_output_mat_60; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_61 = Calc8x8_io_output_mat_61; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_62 = Calc8x8_io_output_mat_62; // @[top.scala 69:26]
  assign Accumu_io_in_from_calc8x8_mat_63 = Calc8x8_io_output_mat_63; // @[top.scala 69:26]
  assign Accumu_io_csum = {{6'd0}, _GEN_152}; // @[Conditional.scala 40:58 para.scala 92:17 top.scala 72:15]
  assign Accumu_io_bias_end_addr = {{6'd0}, _GEN_152}; // @[Conditional.scala 40:58 para.scala 92:17 top.scala 72:15]
  assign Accumu_io_bias_in = ROMBias_io_out; // @[top.scala 76:18]
  assign Accumu_io_is_in_use = 3'h0 == state; // @[Conditional.scala 37:30]
  assign Quant_clock = clock;
  assign Quant_reset = reset;
  assign Quant_io_valid_in = Accumu_io_valid_out; // @[top.scala 81:20]
  assign Quant_io_flag_job = 3'h0 == state; // @[Conditional.scala 37:30]
  assign Quant_io_in_from_accumu_mat_0 = Accumu_io_result_mat_0; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_1 = Accumu_io_result_mat_1; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_2 = Accumu_io_result_mat_2; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_3 = Accumu_io_result_mat_3; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_4 = Accumu_io_result_mat_4; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_5 = Accumu_io_result_mat_5; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_6 = Accumu_io_result_mat_6; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_7 = Accumu_io_result_mat_7; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_8 = Accumu_io_result_mat_8; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_9 = Accumu_io_result_mat_9; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_10 = Accumu_io_result_mat_10; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_11 = Accumu_io_result_mat_11; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_12 = Accumu_io_result_mat_12; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_13 = Accumu_io_result_mat_13; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_14 = Accumu_io_result_mat_14; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_15 = Accumu_io_result_mat_15; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_16 = Accumu_io_result_mat_16; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_17 = Accumu_io_result_mat_17; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_18 = Accumu_io_result_mat_18; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_19 = Accumu_io_result_mat_19; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_20 = Accumu_io_result_mat_20; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_21 = Accumu_io_result_mat_21; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_22 = Accumu_io_result_mat_22; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_23 = Accumu_io_result_mat_23; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_24 = Accumu_io_result_mat_24; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_25 = Accumu_io_result_mat_25; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_26 = Accumu_io_result_mat_26; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_27 = Accumu_io_result_mat_27; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_28 = Accumu_io_result_mat_28; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_29 = Accumu_io_result_mat_29; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_30 = Accumu_io_result_mat_30; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_31 = Accumu_io_result_mat_31; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_32 = Accumu_io_result_mat_32; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_33 = Accumu_io_result_mat_33; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_34 = Accumu_io_result_mat_34; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_35 = Accumu_io_result_mat_35; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_36 = Accumu_io_result_mat_36; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_37 = Accumu_io_result_mat_37; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_38 = Accumu_io_result_mat_38; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_39 = Accumu_io_result_mat_39; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_40 = Accumu_io_result_mat_40; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_41 = Accumu_io_result_mat_41; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_42 = Accumu_io_result_mat_42; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_43 = Accumu_io_result_mat_43; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_44 = Accumu_io_result_mat_44; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_45 = Accumu_io_result_mat_45; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_46 = Accumu_io_result_mat_46; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_47 = Accumu_io_result_mat_47; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_48 = Accumu_io_result_mat_48; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_49 = Accumu_io_result_mat_49; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_50 = Accumu_io_result_mat_50; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_51 = Accumu_io_result_mat_51; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_52 = Accumu_io_result_mat_52; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_53 = Accumu_io_result_mat_53; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_54 = Accumu_io_result_mat_54; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_55 = Accumu_io_result_mat_55; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_56 = Accumu_io_result_mat_56; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_57 = Accumu_io_result_mat_57; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_58 = Accumu_io_result_mat_58; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_59 = Accumu_io_result_mat_59; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_60 = Accumu_io_result_mat_60; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_61 = Accumu_io_result_mat_61; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_62 = Accumu_io_result_mat_62; // @[top.scala 80:26]
  assign Quant_io_in_from_accumu_mat_63 = Accumu_io_result_mat_63; // @[top.scala 80:26]
  assign Quant_io_quant_in_in_q = _T ? 6'h10 : 6'h0; // @[Conditional.scala 40:58 para.scala 102:25 top.scala 83:20]
  assign Quant_io_quant_in_out_q = _T ? 6'h10 : 6'h0; // @[Conditional.scala 40:58 para.scala 103:26 top.scala 83:20]
  assign WriteSwitch_io_valid_in_0 = Quant_io_valid_out; // @[top.scala 97:30]
  assign WriteSwitch_io_input_0_mat_0 = Quant_io_result_mat_0; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_1 = Quant_io_result_mat_1; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_2 = Quant_io_result_mat_2; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_3 = Quant_io_result_mat_3; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_4 = Quant_io_result_mat_4; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_5 = Quant_io_result_mat_5; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_6 = Quant_io_result_mat_6; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_7 = Quant_io_result_mat_7; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_8 = Quant_io_result_mat_8; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_9 = Quant_io_result_mat_9; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_10 = Quant_io_result_mat_10; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_11 = Quant_io_result_mat_11; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_12 = Quant_io_result_mat_12; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_13 = Quant_io_result_mat_13; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_14 = Quant_io_result_mat_14; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_15 = Quant_io_result_mat_15; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_16 = Quant_io_result_mat_16; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_17 = Quant_io_result_mat_17; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_18 = Quant_io_result_mat_18; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_19 = Quant_io_result_mat_19; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_20 = Quant_io_result_mat_20; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_21 = Quant_io_result_mat_21; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_22 = Quant_io_result_mat_22; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_23 = Quant_io_result_mat_23; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_24 = Quant_io_result_mat_24; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_25 = Quant_io_result_mat_25; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_26 = Quant_io_result_mat_26; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_27 = Quant_io_result_mat_27; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_28 = Quant_io_result_mat_28; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_29 = Quant_io_result_mat_29; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_30 = Quant_io_result_mat_30; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_31 = Quant_io_result_mat_31; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_32 = Quant_io_result_mat_32; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_33 = Quant_io_result_mat_33; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_34 = Quant_io_result_mat_34; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_35 = Quant_io_result_mat_35; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_36 = Quant_io_result_mat_36; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_37 = Quant_io_result_mat_37; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_38 = Quant_io_result_mat_38; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_39 = Quant_io_result_mat_39; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_40 = Quant_io_result_mat_40; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_41 = Quant_io_result_mat_41; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_42 = Quant_io_result_mat_42; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_43 = Quant_io_result_mat_43; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_44 = Quant_io_result_mat_44; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_45 = Quant_io_result_mat_45; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_46 = Quant_io_result_mat_46; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_47 = Quant_io_result_mat_47; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_48 = Quant_io_result_mat_48; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_49 = Quant_io_result_mat_49; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_50 = Quant_io_result_mat_50; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_51 = Quant_io_result_mat_51; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_52 = Quant_io_result_mat_52; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_53 = Quant_io_result_mat_53; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_54 = Quant_io_result_mat_54; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_55 = Quant_io_result_mat_55; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_56 = Quant_io_result_mat_56; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_57 = Quant_io_result_mat_57; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_58 = Quant_io_result_mat_58; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_59 = Quant_io_result_mat_59; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_60 = Quant_io_result_mat_60; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_61 = Quant_io_result_mat_61; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_62 = Quant_io_result_mat_62; // @[top.scala 104:27]
  assign WriteSwitch_io_input_0_mat_63 = Quant_io_result_mat_63; // @[top.scala 104:27]
  assign RealWriter_clock = clock;
  assign RealWriter_reset = reset;
  assign RealWriter_io_valid_in = WriteSwitch_io_valid_out; // @[top.scala 109:21]
  assign RealWriter_io_flag_job = 3'h0 == state; // @[Conditional.scala 37:30]
  assign RealWriter_io_in_from_quant_mat_0 = WriteSwitch_io_output_mat_0; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_1 = WriteSwitch_io_output_mat_1; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_2 = WriteSwitch_io_output_mat_2; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_3 = WriteSwitch_io_output_mat_3; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_4 = WriteSwitch_io_output_mat_4; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_5 = WriteSwitch_io_output_mat_5; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_6 = WriteSwitch_io_output_mat_6; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_7 = WriteSwitch_io_output_mat_7; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_8 = WriteSwitch_io_output_mat_8; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_9 = WriteSwitch_io_output_mat_9; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_10 = WriteSwitch_io_output_mat_10; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_11 = WriteSwitch_io_output_mat_11; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_12 = WriteSwitch_io_output_mat_12; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_13 = WriteSwitch_io_output_mat_13; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_14 = WriteSwitch_io_output_mat_14; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_15 = WriteSwitch_io_output_mat_15; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_16 = WriteSwitch_io_output_mat_16; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_17 = WriteSwitch_io_output_mat_17; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_18 = WriteSwitch_io_output_mat_18; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_19 = WriteSwitch_io_output_mat_19; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_20 = WriteSwitch_io_output_mat_20; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_21 = WriteSwitch_io_output_mat_21; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_22 = WriteSwitch_io_output_mat_22; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_23 = WriteSwitch_io_output_mat_23; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_24 = WriteSwitch_io_output_mat_24; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_25 = WriteSwitch_io_output_mat_25; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_26 = WriteSwitch_io_output_mat_26; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_27 = WriteSwitch_io_output_mat_27; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_28 = WriteSwitch_io_output_mat_28; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_29 = WriteSwitch_io_output_mat_29; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_30 = WriteSwitch_io_output_mat_30; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_31 = WriteSwitch_io_output_mat_31; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_32 = WriteSwitch_io_output_mat_32; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_33 = WriteSwitch_io_output_mat_33; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_34 = WriteSwitch_io_output_mat_34; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_35 = WriteSwitch_io_output_mat_35; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_36 = WriteSwitch_io_output_mat_36; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_37 = WriteSwitch_io_output_mat_37; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_38 = WriteSwitch_io_output_mat_38; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_39 = WriteSwitch_io_output_mat_39; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_40 = WriteSwitch_io_output_mat_40; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_41 = WriteSwitch_io_output_mat_41; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_42 = WriteSwitch_io_output_mat_42; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_43 = WriteSwitch_io_output_mat_43; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_44 = WriteSwitch_io_output_mat_44; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_45 = WriteSwitch_io_output_mat_45; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_46 = WriteSwitch_io_output_mat_46; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_47 = WriteSwitch_io_output_mat_47; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_48 = WriteSwitch_io_output_mat_48; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_49 = WriteSwitch_io_output_mat_49; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_50 = WriteSwitch_io_output_mat_50; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_51 = WriteSwitch_io_output_mat_51; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_52 = WriteSwitch_io_output_mat_52; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_53 = WriteSwitch_io_output_mat_53; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_54 = WriteSwitch_io_output_mat_54; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_55 = WriteSwitch_io_output_mat_55; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_56 = WriteSwitch_io_output_mat_56; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_57 = WriteSwitch_io_output_mat_57; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_58 = WriteSwitch_io_output_mat_58; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_59 = WriteSwitch_io_output_mat_59; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_60 = WriteSwitch_io_output_mat_60; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_61 = WriteSwitch_io_output_mat_61; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_62 = WriteSwitch_io_output_mat_62; // @[top.scala 108:26]
  assign RealWriter_io_in_from_quant_mat_63 = WriteSwitch_io_output_mat_63; // @[top.scala 108:26]
  assign RealWriter_io_job_job_0_big_begin_addr = _T ? 10'h40 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_big_max_addr = _T ? 10'h383 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_big_cnt_ic_end = _T ? 10'hf : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_big_a = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_0_begin_addr = _T ? 10'h20 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_0_max_addr = _T ? 10'h1c1 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_0_cnt_y_end = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_0_cnt_ic_end = _T ? 10'hf : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_0_a = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_0_ano_bank_id = _T ? 3'h2 : 3'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_1_begin_addr = _T ? 10'h20 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_1_max_addr = _T ? 10'h1c1 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_1_bank_id = _T ? 3'h1 : 3'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_1_cnt_y_end = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_1_cnt_ic_end = _T ? 10'hf : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_1_a = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_0_small_1_ano_bank_id = _T ? 3'h3 : 3'h0; // @[Conditional.scala 40:58 para.scala 114:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_big_begin_addr = _T ? 10'h40 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_big_max_addr = _T ? 10'h383 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_big_bank_id = _T ? 3'h1 : 3'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_big_cnt_ic_end = _T ? 10'hf : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_big_a = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_0_begin_addr = _T ? 10'h20 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_0_max_addr = _T ? 10'h1c1 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_0_bank_id = _T ? 3'h4 : 3'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_0_cnt_y_end = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_0_cnt_ic_end = _T ? 10'hf : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_0_a = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_0_ano_bank_id = _T ? 3'h6 : 3'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_1_begin_addr = _T ? 10'h20 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_1_max_addr = _T ? 10'h1c1 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_1_bank_id = _T ? 3'h5 : 3'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_1_cnt_y_end = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_1_cnt_ic_end = _T ? 10'hf : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_1_a = _T ? 10'h1 : 10'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_job_1_small_1_ano_bank_id = _T ? 3'h7 : 3'h0; // @[Conditional.scala 40:58 para.scala 121:23 top.scala 111:16]
  assign RealWriter_io_job_out_chan = _T ? 10'h10 : 10'h0; // @[Conditional.scala 40:58 para.scala 128:25 top.scala 111:16]
  assign ROMWeight_clock = clock;
  assign ROMWeight_io_addr = WeightReader_io_addr; // @[top.scala 47:21]
  assign ROMBias_clock = clock;
  assign ROMBias_io_addr = Accumu_io_bias_addr[7:0]; // @[top.scala 75:19]
  assign RAMGroup_clock = clock;
  assign RAMGroup_reset = reset;
  assign RAMGroup_io_rd_valid_in = GraphReader_1_io_valid_out; // @[top.scala 37:22]
  assign RAMGroup_io_rd_addr1_addrs_0_bank_id = GraphReader_io_to_banks_addrs_0_bank_id; // @[top.scala 31:19]
  assign RAMGroup_io_rd_addr1_addrs_1_addr = GraphReader_io_to_banks_addrs_1_addr; // @[top.scala 31:19]
  assign RAMGroup_io_rd_addr2_addrs_1_addr = GraphReader_1_io_to_banks_addrs_1_addr; // @[top.scala 38:19]
  always @(posedge clock) begin
    if (reset) begin // @[top.scala 134:26]
      counter_ccnt <= 10'h0; // @[top.scala 134:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      counter_ccnt <= 10'h0; // @[utils.scala 23:14]
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (RealWriter_io_valid_out) begin // @[top.scala 152:35]
        counter_ccnt <= _counter_ccnt_T_2; // @[utils.scala 18:14]
      end
    end
    if (reset) begin // @[top.scala 134:26]
      counter_cend <= 10'h0; // @[top.scala 134:26]
    end else if (_T) begin // @[Conditional.scala 40:58]
      counter_cend <= 10'h3f; // @[utils.scala 22:14]
    end
    if (reset) begin // @[top.scala 135:24]
      state <= 3'h0; // @[top.scala 135:24]
    end else if (_T) begin // @[Conditional.scala 40:58]
      state <= 3'h1; // @[top.scala 149:19]
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (RealWriter_io_valid_out) begin // @[top.scala 152:35]
        state <= _GEN_0;
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      state <= 3'h2; // @[top.scala 164:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter_ccnt = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  counter_cend = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
